module tt_um_sky130_as_sc_hs_dyn_test (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net21;
 wire net22;
 wire net23;

 sky130_as_sc_hs__xnor2_2 _35_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(uio_out[4]),
    .Y(_16_),
    .B(uio_out[2]));
 sky130_as_sc_hs__xnor2_2 _36_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(uio_out[5]),
    .Y(_17_),
    .B(uio_out[7]));
 sky130_as_sc_hs__xnor2_2 _37_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_16_),
    .Y(_18_),
    .B(_17_));
 sky130_as_sc_hs__nor2_2 _38_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net2),
    .B(net12),
    .Y(_19_));
 sky130_as_sc_hs__aoi21_2 _39_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net11),
    .B(_18_),
    .C(_19_),
    .Y(_00_));
 sky130_as_sc_hs__mux2_2 _40_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net12),
    .B(uo_out[0]),
    .A(net3),
    .Y(_20_));
 sky130_as_sc_hs__buff_2 _41_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_20_),
    .Y(_01_));
 sky130_as_sc_hs__mux2_2 _42_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net12),
    .B(uo_out[1]),
    .A(net4),
    .Y(_21_));
 sky130_as_sc_hs__buff_2 _43_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_21_),
    .Y(_02_));
 sky130_as_sc_hs__mux2_2 _44_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net12),
    .B(uo_out[2]),
    .A(net5),
    .Y(_22_));
 sky130_as_sc_hs__buff_2 _45_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_22_),
    .Y(_03_));
 sky130_as_sc_hs__mux2_2 _46_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net12),
    .B(uo_out[3]),
    .A(net6),
    .Y(_23_));
 sky130_as_sc_hs__buff_2 _47_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_23_),
    .Y(_04_));
 sky130_as_sc_hs__mux2_2 _48_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net1),
    .B(uo_out[4]),
    .A(net7),
    .Y(_24_));
 sky130_as_sc_hs__buff_2 _49_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_24_),
    .Y(_05_));
 sky130_as_sc_hs__mux2_2 _50_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net1),
    .B(uo_out[5]),
    .A(net8),
    .Y(_25_));
 sky130_as_sc_hs__buff_2 _51_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_25_),
    .Y(_06_));
 sky130_as_sc_hs__mux2_2 _52_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net11),
    .B(uo_out[6]),
    .A(net9),
    .Y(_26_));
 sky130_as_sc_hs__buff_2 _53_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_26_),
    .Y(_07_));
 sky130_as_sc_hs__nand2b_2 _54_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(net11),
    .Y(_27_),
    .A(uo_out[7]));
 sky130_as_sc_hs__buff_2 _55_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_27_),
    .Y(_08_));
 sky130_as_sc_hs__and2_2 _56_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net10),
    .B(uio_out[0]),
    .Y(_28_));
 sky130_as_sc_hs__buff_2 _57_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_28_),
    .Y(_09_));
 sky130_as_sc_hs__and2_2 _58_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net10),
    .B(uio_out[1]),
    .Y(_29_));
 sky130_as_sc_hs__buff_2 _59_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_29_),
    .Y(_10_));
 sky130_as_sc_hs__and2_2 _60_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net21),
    .B(net10),
    .Y(_30_));
 sky130_as_sc_hs__buff_2 _61_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_30_),
    .Y(_11_));
 sky130_as_sc_hs__and2_2 _62_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net10),
    .B(uio_out[3]),
    .Y(_31_));
 sky130_as_sc_hs__buff_2 _63_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_31_),
    .Y(_12_));
 sky130_as_sc_hs__and2_2 _64_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net22),
    .B(net10),
    .Y(_32_));
 sky130_as_sc_hs__buff_2 _65_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_32_),
    .Y(_13_));
 sky130_as_sc_hs__and2_2 _66_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net23),
    .B(net10),
    .Y(_33_));
 sky130_as_sc_hs__buff_2 _67_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_33_),
    .Y(_14_));
 sky130_as_sc_hs__and2_2 _68_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net10),
    .B(uio_out[6]),
    .Y(_34_));
 sky130_as_sc_hs__buff_2 _69_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_34_),
    .Y(_15_));
 sky130_as_sc_hs__dyn_dfxtp_4 _70_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_0__leaf_clk),
    .D(_08_),
    .Q(uio_out[0]));
 sky130_as_sc_hs__dyn_dfxtp_4 _71_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_0__leaf_clk),
    .D(_09_),
    .Q(uio_out[1]));
 sky130_as_sc_hs__dyn_dfxtp_4 _72_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_0__leaf_clk),
    .D(_10_),
    .Q(uio_out[2]));
 sky130_as_sc_hs__dyn_dfxtp_4 _73_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_0__leaf_clk),
    .D(_11_),
    .Q(uio_out[3]));
 sky130_as_sc_hs__dyn_dfxtp_4 _74_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_0__leaf_clk),
    .D(_12_),
    .Q(uio_out[4]));
 sky130_as_sc_hs__dyn_dfxtp_4 _75_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_0__leaf_clk),
    .D(_13_),
    .Q(uio_out[5]));
 sky130_as_sc_hs__dyn_dfxtp_4 _76_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_0__leaf_clk),
    .D(_14_),
    .Q(uio_out[6]));
 sky130_as_sc_hs__dyn_dfxtp_4 _77_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_0__leaf_clk),
    .D(_15_),
    .Q(uio_out[7]));
 sky130_as_sc_hs__dyn_dfxtp_4 _78_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_1__leaf_clk),
    .D(_00_),
    .Q(uo_out[0]));
 sky130_as_sc_hs__dyn_dfxtp_4 _79_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_1__leaf_clk),
    .D(_01_),
    .Q(uo_out[1]));
 sky130_as_sc_hs__dyn_dfxtp_4 _80_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_1__leaf_clk),
    .D(_02_),
    .Q(uo_out[2]));
 sky130_as_sc_hs__dyn_dfxtp_4 _81_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_1__leaf_clk),
    .D(_03_),
    .Q(uo_out[3]));
 sky130_as_sc_hs__dyn_dfxtp_4 _82_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_1__leaf_clk),
    .D(_04_),
    .Q(uo_out[4]));
 sky130_as_sc_hs__dyn_dfxtp_4 _83_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_1__leaf_clk),
    .D(_05_),
    .Q(uo_out[5]));
 sky130_as_sc_hs__dyn_dfxtp_4 _84_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_1__leaf_clk),
    .D(_06_),
    .Q(uo_out[6]));
 sky130_as_sc_hs__dyn_dfxtp_4 _85_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_1_1__leaf_clk),
    .D(_07_),
    .Q(uo_out[7]));
 sky130_as_sc_hs__tieh tt_um_sky130_as_sc_hs_dyn_test_14 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ONE(net14));
 sky130_as_sc_hs__tieh tt_um_sky130_as_sc_hs_dyn_test_15 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ONE(net15));
 sky130_as_sc_hs__tieh tt_um_sky130_as_sc_hs_dyn_test_16 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ONE(net16));
 sky130_as_sc_hs__tieh tt_um_sky130_as_sc_hs_dyn_test_17 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ONE(net17));
 sky130_as_sc_hs__tieh tt_um_sky130_as_sc_hs_dyn_test_18 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ONE(net18));
 sky130_as_sc_hs__tieh tt_um_sky130_as_sc_hs_dyn_test_19 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ONE(net19));
 sky130_as_sc_hs__tieh tt_um_sky130_as_sc_hs_dyn_test_20 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ONE(net20));
 sky130_as_sc_hs__clkbuff_11 clkbuf_0_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clk),
    .Y(clknet_0_clk));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_0_Right_0 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_1_Right_1 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_2_Right_2 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_3_Right_3 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_4_Right_4 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_5_Right_5 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_6_Right_6 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_7_Right_7 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_8_Right_8 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_9_Right_9 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_10_Right_10 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_11_Right_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_12_Right_12 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_13_Right_13 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_14_Right_14 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_15_Right_15 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_16_Right_16 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_17_Right_17 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_18_Right_18 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_19_Right_19 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_20_Right_20 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_21_Right_21 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_22_Right_22 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_23_Right_23 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_24_Right_24 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_25_Right_25 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_26_Right_26 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_27_Right_27 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_28_Right_28 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_29_Right_29 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_30_Right_30 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_31_Right_31 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_32_Right_32 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_33_Right_33 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_34_Right_34 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_35_Right_35 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_36_Right_36 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_37_Right_37 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_38_Right_38 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_0_Left_39 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_1_Left_40 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_2_Left_41 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_3_Left_42 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_4_Left_43 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_5_Left_44 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_6_Left_45 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_7_Left_46 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_8_Left_47 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_9_Left_48 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_10_Left_49 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_11_Left_50 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_12_Left_51 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_13_Left_52 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_14_Left_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_15_Left_54 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_16_Left_55 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_17_Left_56 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_18_Left_57 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_19_Left_58 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_20_Left_59 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_21_Left_60 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_22_Left_61 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_23_Left_62 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_24_Left_63 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_25_Left_64 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_26_Left_65 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_27_Left_66 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_28_Left_67 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_29_Left_68 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_30_Left_69 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_31_Left_70 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_32_Left_71 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_33_Left_72 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_34_Left_73 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_35_Left_74 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_36_Left_75 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_37_Left_76 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_38_Left_77 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_78 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_79 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_80 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_81 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_82 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_83 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_84 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_85 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_86 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_87 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_88 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_89 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_90 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_91 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_92 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_93 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_94 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_95 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_96 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_97 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_98 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_99 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_100 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_101 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_102 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_103 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_104 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_105 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_106 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_107 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_108 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_109 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_110 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_111 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_112 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_113 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_114 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_115 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_116 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_117 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_118 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_119 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_120 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_121 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_122 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_123 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_124 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_125 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_126 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_127 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_128 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_129 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_130 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_131 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_132 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_133 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_134 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_135 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_136 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_137 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_138 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_139 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_140 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_141 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_142 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_143 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_144 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_145 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_146 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_147 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_148 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_149 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_150 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_151 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_152 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_153 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_154 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_155 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_156 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_157 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_158 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_159 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_160 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_161 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_162 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_163 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_164 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_165 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_166 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_167 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_168 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_169 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_170 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_171 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_172 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_173 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_174 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_175 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_176 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_177 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_178 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_179 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_180 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_181 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_182 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_183 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_184 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_185 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_186 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_187 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_188 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_189 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_190 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_191 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_192 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_193 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_194 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_195 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_196 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_197 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_198 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_199 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_200 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_201 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_202 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_203 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_204 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_205 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_206 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_207 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_208 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_209 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_210 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_211 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_212 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_213 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_214 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_215 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_216 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_217 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_218 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_219 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_220 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_221 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_222 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_223 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_224 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_225 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_226 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_227 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_228 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_229 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_230 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_231 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_232 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_233 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_234 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_235 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_236 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_237 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_238 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_239 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_240 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_241 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_242 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_243 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_244 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_245 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_246 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_247 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_248 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_249 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_250 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_251 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_252 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_253 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_254 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_255 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_256 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_257 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_258 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_259 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_260 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_261 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_262 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_263 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_264 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_265 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_266 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_267 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_268 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_269 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_270 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_271 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_272 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_273 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_274 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_275 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_276 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_277 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_278 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_279 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_280 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_281 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_282 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_283 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_284 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_285 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_286 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_287 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_288 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_289 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_290 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_291 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_292 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_293 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_294 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_295 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_296 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_297 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_298 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_299 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_300 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_301 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_302 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__buff_2 input1 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(rst_n),
    .Y(net1));
 sky130_as_sc_hs__buff_2 input2 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[0]),
    .Y(net2));
 sky130_as_sc_hs__buff_2 input3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[1]),
    .Y(net3));
 sky130_as_sc_hs__buff_2 input4 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[2]),
    .Y(net4));
 sky130_as_sc_hs__buff_2 input5 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[3]),
    .Y(net5));
 sky130_as_sc_hs__buff_2 input6 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[4]),
    .Y(net6));
 sky130_as_sc_hs__buff_2 input7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[5]),
    .Y(net7));
 sky130_as_sc_hs__buff_2 input8 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[6]),
    .Y(net8));
 sky130_as_sc_hs__buff_2 input9 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[7]),
    .Y(net9));
 sky130_as_sc_hs__buff_2 fanout10 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net12),
    .Y(net10));
 sky130_as_sc_hs__buff_2 fanout11 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net12),
    .Y(net11));
 sky130_as_sc_hs__buff_4 fanout12 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net1),
    .Y(net12));
 sky130_as_sc_hs__tieh tt_um_sky130_as_sc_hs_dyn_test_13 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ONE(net13));
 sky130_as_sc_hs__clkbuff_11 clkbuf_1_0__f_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_0_clk),
    .Y(clknet_1_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_11 clkbuf_1_1__f_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_0_clk),
    .Y(clknet_1_1__leaf_clk));
 sky130_as_sc_hs__buff_2 hold1 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_out[2]),
    .Y(net21));
 sky130_as_sc_hs__buff_2 hold2 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_out[4]),
    .Y(net22));
 sky130_as_sc_hs__buff_2 hold3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_out[5]),
    .Y(net23));
 sky130_as_sc_hs__decap_16 FILLER_0_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_0_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_0_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_45 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_73 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_129 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_157 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_185 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_213 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_269 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_297 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_0_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_1_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_1_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_2_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_2_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_2_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_2_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_3_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_3_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_4_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_4_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_4_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_4_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_5_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_5_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_6_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_6_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_6_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_6_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_7_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_7_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_8_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_8_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_8_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_8_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_9_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_9_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_10_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_10_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_10_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_10_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_11_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_11_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_11_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_11_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_11_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_11_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_12_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_12_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_12_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_12_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_13_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_13_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_14_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_14_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_14_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_14_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_14_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_14_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_14_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_14_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_14_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_15_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_15_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_15_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_15_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_15_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_15_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_16_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_16_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_16_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_16_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_16_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_16_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_16_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_16_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_16_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_17_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_17_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_17_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_17_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_17_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_17_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_17_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_17_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_17_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_18_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_18_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_18_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_18_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_18_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_18_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_18_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_18_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_18_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_19_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_19_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_19_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_19_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_19_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_19_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_20_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_20_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_20_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_20_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_20_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_20_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_20_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_20_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_20_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_21_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_21_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_21_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_21_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_21_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_22_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_22_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_22_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_22_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_22_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_22_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_22_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_22_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_22_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_23_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_23_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_23_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_23_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_23_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_23_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_24_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_24_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_24_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_24_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_24_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_24_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_24_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_24_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_24_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_25_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_25_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_25_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_25_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_25_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_26_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_26_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_26_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_26_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_26_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_26_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_26_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_26_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_26_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_27_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_27_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_27_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_27_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_27_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_27_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_27_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_27_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_27_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_28_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_28_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_28_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_28_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_28_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_28_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_28_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_28_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_28_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_29_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_29_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_29_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_29_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_29_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_30_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_30_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_30_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_30_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_30_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_30_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_30_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_30_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_30_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_31_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_31_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_31_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_31_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_31_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_31_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_32_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_32_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_32_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_32_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_32_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_32_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_32_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_32_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_32_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_33_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_33_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_33_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_33_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_33_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_33_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_34_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_34_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_34_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_117 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_34_132 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_34_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_34_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_34_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_34_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_34_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_35_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_35_89 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_97 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_35_101 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_35_146 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_35_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_35_185 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_193 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_35_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_35_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_35_245 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_35_268 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_276 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_35_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_36_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_36_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_36_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_156 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_176 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_36_194 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_240 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_276 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_292 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_36_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_36_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_173 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_37_229 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_37_278 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_300 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_316 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_332 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_38_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_38_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_38_45 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_38_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_64 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_38_70 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_38_76 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_38_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_88 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_135 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_146 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_38_155 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_185 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_38_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_223 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_251 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_278 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_38_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
endmodule
