module tt_um_sky130_as_sc_hs (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \A[0] ;
 wire \A[1] ;
 wire \A[2] ;
 wire \A[3] ;
 wire \A[4] ;
 wire \A[5] ;
 wire \B[0] ;
 wire \B[1] ;
 wire \B[2] ;
 wire \B[3] ;
 wire \B[4] ;
 wire \B[5] ;
 wire CS_ROM;
 wire HCF;
 wire \MAR[0] ;
 wire \MAR[1] ;
 wire \MAR[2] ;
 wire \MAR[3] ;
 wire \MAR[4] ;
 wire \MAR[5] ;
 wire \PC[0] ;
 wire \PC[10] ;
 wire \PC[11] ;
 wire \PC[1] ;
 wire \PC[2] ;
 wire \PC[3] ;
 wire \PC[4] ;
 wire \PC[5] ;
 wire \PC[6] ;
 wire \PC[7] ;
 wire \PC[8] ;
 wire \PC[9] ;
 wire \P[0] ;
 wire \P[1] ;
 wire \P[2] ;
 wire \P[3] ;
 wire \P[4] ;
 wire \P[5] ;
 wire \RAM[0][0] ;
 wire \RAM[0][1] ;
 wire \RAM[0][2] ;
 wire \RAM[0][3] ;
 wire \RAM[0][4] ;
 wire \RAM[0][5] ;
 wire \RAM[10][0] ;
 wire \RAM[10][1] ;
 wire \RAM[10][2] ;
 wire \RAM[10][3] ;
 wire \RAM[10][4] ;
 wire \RAM[10][5] ;
 wire \RAM[11][0] ;
 wire \RAM[11][1] ;
 wire \RAM[11][2] ;
 wire \RAM[11][3] ;
 wire \RAM[11][4] ;
 wire \RAM[11][5] ;
 wire \RAM[12][0] ;
 wire \RAM[12][1] ;
 wire \RAM[12][2] ;
 wire \RAM[12][3] ;
 wire \RAM[12][4] ;
 wire \RAM[12][5] ;
 wire \RAM[13][0] ;
 wire \RAM[13][1] ;
 wire \RAM[13][2] ;
 wire \RAM[13][3] ;
 wire \RAM[13][4] ;
 wire \RAM[13][5] ;
 wire \RAM[14][0] ;
 wire \RAM[14][1] ;
 wire \RAM[14][2] ;
 wire \RAM[14][3] ;
 wire \RAM[14][4] ;
 wire \RAM[14][5] ;
 wire \RAM[15][0] ;
 wire \RAM[15][1] ;
 wire \RAM[15][2] ;
 wire \RAM[15][3] ;
 wire \RAM[15][4] ;
 wire \RAM[15][5] ;
 wire \RAM[16][0] ;
 wire \RAM[16][1] ;
 wire \RAM[16][2] ;
 wire \RAM[16][3] ;
 wire \RAM[16][4] ;
 wire \RAM[16][5] ;
 wire \RAM[17][0] ;
 wire \RAM[17][1] ;
 wire \RAM[17][2] ;
 wire \RAM[17][3] ;
 wire \RAM[17][4] ;
 wire \RAM[17][5] ;
 wire \RAM[18][0] ;
 wire \RAM[18][1] ;
 wire \RAM[18][2] ;
 wire \RAM[18][3] ;
 wire \RAM[18][4] ;
 wire \RAM[18][5] ;
 wire \RAM[19][0] ;
 wire \RAM[19][1] ;
 wire \RAM[19][2] ;
 wire \RAM[19][3] ;
 wire \RAM[19][4] ;
 wire \RAM[19][5] ;
 wire \RAM[1][0] ;
 wire \RAM[1][1] ;
 wire \RAM[1][2] ;
 wire \RAM[1][3] ;
 wire \RAM[1][4] ;
 wire \RAM[1][5] ;
 wire \RAM[20][0] ;
 wire \RAM[20][1] ;
 wire \RAM[20][2] ;
 wire \RAM[20][3] ;
 wire \RAM[20][4] ;
 wire \RAM[20][5] ;
 wire \RAM[21][0] ;
 wire \RAM[21][1] ;
 wire \RAM[21][2] ;
 wire \RAM[21][3] ;
 wire \RAM[21][4] ;
 wire \RAM[21][5] ;
 wire \RAM[22][0] ;
 wire \RAM[22][1] ;
 wire \RAM[22][2] ;
 wire \RAM[22][3] ;
 wire \RAM[22][4] ;
 wire \RAM[22][5] ;
 wire \RAM[23][0] ;
 wire \RAM[23][1] ;
 wire \RAM[23][2] ;
 wire \RAM[23][3] ;
 wire \RAM[23][4] ;
 wire \RAM[23][5] ;
 wire \RAM[24][0] ;
 wire \RAM[24][1] ;
 wire \RAM[24][2] ;
 wire \RAM[24][3] ;
 wire \RAM[24][4] ;
 wire \RAM[24][5] ;
 wire \RAM[25][0] ;
 wire \RAM[25][1] ;
 wire \RAM[25][2] ;
 wire \RAM[25][3] ;
 wire \RAM[25][4] ;
 wire \RAM[25][5] ;
 wire \RAM[26][0] ;
 wire \RAM[26][1] ;
 wire \RAM[26][2] ;
 wire \RAM[26][3] ;
 wire \RAM[26][4] ;
 wire \RAM[26][5] ;
 wire \RAM[27][0] ;
 wire \RAM[27][1] ;
 wire \RAM[27][2] ;
 wire \RAM[27][3] ;
 wire \RAM[27][4] ;
 wire \RAM[27][5] ;
 wire \RAM[28][0] ;
 wire \RAM[28][1] ;
 wire \RAM[28][2] ;
 wire \RAM[28][3] ;
 wire \RAM[28][4] ;
 wire \RAM[28][5] ;
 wire \RAM[29][0] ;
 wire \RAM[29][1] ;
 wire \RAM[29][2] ;
 wire \RAM[29][3] ;
 wire \RAM[29][4] ;
 wire \RAM[29][5] ;
 wire \RAM[2][0] ;
 wire \RAM[2][1] ;
 wire \RAM[2][2] ;
 wire \RAM[2][3] ;
 wire \RAM[2][4] ;
 wire \RAM[2][5] ;
 wire \RAM[30][0] ;
 wire \RAM[30][1] ;
 wire \RAM[30][2] ;
 wire \RAM[30][3] ;
 wire \RAM[30][4] ;
 wire \RAM[30][5] ;
 wire \RAM[31][0] ;
 wire \RAM[31][1] ;
 wire \RAM[31][2] ;
 wire \RAM[31][3] ;
 wire \RAM[31][4] ;
 wire \RAM[31][5] ;
 wire \RAM[32][0] ;
 wire \RAM[32][1] ;
 wire \RAM[32][2] ;
 wire \RAM[32][3] ;
 wire \RAM[32][4] ;
 wire \RAM[32][5] ;
 wire \RAM[33][0] ;
 wire \RAM[33][1] ;
 wire \RAM[33][2] ;
 wire \RAM[33][3] ;
 wire \RAM[33][4] ;
 wire \RAM[33][5] ;
 wire \RAM[34][0] ;
 wire \RAM[34][1] ;
 wire \RAM[34][2] ;
 wire \RAM[34][3] ;
 wire \RAM[34][4] ;
 wire \RAM[34][5] ;
 wire \RAM[35][0] ;
 wire \RAM[35][1] ;
 wire \RAM[35][2] ;
 wire \RAM[35][3] ;
 wire \RAM[35][4] ;
 wire \RAM[35][5] ;
 wire \RAM[36][0] ;
 wire \RAM[36][1] ;
 wire \RAM[36][2] ;
 wire \RAM[36][3] ;
 wire \RAM[36][4] ;
 wire \RAM[36][5] ;
 wire \RAM[37][0] ;
 wire \RAM[37][1] ;
 wire \RAM[37][2] ;
 wire \RAM[37][3] ;
 wire \RAM[37][4] ;
 wire \RAM[37][5] ;
 wire \RAM[38][0] ;
 wire \RAM[38][1] ;
 wire \RAM[38][2] ;
 wire \RAM[38][3] ;
 wire \RAM[38][4] ;
 wire \RAM[38][5] ;
 wire \RAM[39][0] ;
 wire \RAM[39][1] ;
 wire \RAM[39][2] ;
 wire \RAM[39][3] ;
 wire \RAM[39][4] ;
 wire \RAM[39][5] ;
 wire \RAM[3][0] ;
 wire \RAM[3][1] ;
 wire \RAM[3][2] ;
 wire \RAM[3][3] ;
 wire \RAM[3][4] ;
 wire \RAM[3][5] ;
 wire \RAM[40][0] ;
 wire \RAM[40][1] ;
 wire \RAM[40][2] ;
 wire \RAM[40][3] ;
 wire \RAM[40][4] ;
 wire \RAM[40][5] ;
 wire \RAM[41][0] ;
 wire \RAM[41][1] ;
 wire \RAM[41][2] ;
 wire \RAM[41][3] ;
 wire \RAM[41][4] ;
 wire \RAM[41][5] ;
 wire \RAM[42][0] ;
 wire \RAM[42][1] ;
 wire \RAM[42][2] ;
 wire \RAM[42][3] ;
 wire \RAM[42][4] ;
 wire \RAM[42][5] ;
 wire \RAM[43][0] ;
 wire \RAM[43][1] ;
 wire \RAM[43][2] ;
 wire \RAM[43][3] ;
 wire \RAM[43][4] ;
 wire \RAM[43][5] ;
 wire \RAM[44][0] ;
 wire \RAM[44][1] ;
 wire \RAM[44][2] ;
 wire \RAM[44][3] ;
 wire \RAM[44][4] ;
 wire \RAM[44][5] ;
 wire \RAM[45][0] ;
 wire \RAM[45][1] ;
 wire \RAM[45][2] ;
 wire \RAM[45][3] ;
 wire \RAM[45][4] ;
 wire \RAM[45][5] ;
 wire \RAM[46][0] ;
 wire \RAM[46][1] ;
 wire \RAM[46][2] ;
 wire \RAM[46][3] ;
 wire \RAM[46][4] ;
 wire \RAM[46][5] ;
 wire \RAM[47][0] ;
 wire \RAM[47][1] ;
 wire \RAM[47][2] ;
 wire \RAM[47][3] ;
 wire \RAM[47][4] ;
 wire \RAM[47][5] ;
 wire \RAM[48][0] ;
 wire \RAM[48][1] ;
 wire \RAM[48][2] ;
 wire \RAM[48][3] ;
 wire \RAM[48][4] ;
 wire \RAM[48][5] ;
 wire \RAM[49][0] ;
 wire \RAM[49][1] ;
 wire \RAM[49][2] ;
 wire \RAM[49][3] ;
 wire \RAM[49][4] ;
 wire \RAM[49][5] ;
 wire \RAM[4][0] ;
 wire \RAM[4][1] ;
 wire \RAM[4][2] ;
 wire \RAM[4][3] ;
 wire \RAM[4][4] ;
 wire \RAM[4][5] ;
 wire \RAM[50][0] ;
 wire \RAM[50][1] ;
 wire \RAM[50][2] ;
 wire \RAM[50][3] ;
 wire \RAM[50][4] ;
 wire \RAM[50][5] ;
 wire \RAM[51][0] ;
 wire \RAM[51][1] ;
 wire \RAM[51][2] ;
 wire \RAM[51][3] ;
 wire \RAM[51][4] ;
 wire \RAM[51][5] ;
 wire \RAM[52][0] ;
 wire \RAM[52][1] ;
 wire \RAM[52][2] ;
 wire \RAM[52][3] ;
 wire \RAM[52][4] ;
 wire \RAM[52][5] ;
 wire \RAM[53][0] ;
 wire \RAM[53][1] ;
 wire \RAM[53][2] ;
 wire \RAM[53][3] ;
 wire \RAM[53][4] ;
 wire \RAM[53][5] ;
 wire \RAM[54][0] ;
 wire \RAM[54][1] ;
 wire \RAM[54][2] ;
 wire \RAM[54][3] ;
 wire \RAM[54][4] ;
 wire \RAM[54][5] ;
 wire \RAM[55][0] ;
 wire \RAM[55][1] ;
 wire \RAM[55][2] ;
 wire \RAM[55][3] ;
 wire \RAM[55][4] ;
 wire \RAM[55][5] ;
 wire \RAM[56][0] ;
 wire \RAM[56][1] ;
 wire \RAM[56][2] ;
 wire \RAM[56][3] ;
 wire \RAM[56][4] ;
 wire \RAM[56][5] ;
 wire \RAM[57][0] ;
 wire \RAM[57][1] ;
 wire \RAM[57][2] ;
 wire \RAM[57][3] ;
 wire \RAM[57][4] ;
 wire \RAM[57][5] ;
 wire \RAM[58][0] ;
 wire \RAM[58][1] ;
 wire \RAM[58][2] ;
 wire \RAM[58][3] ;
 wire \RAM[58][4] ;
 wire \RAM[58][5] ;
 wire \RAM[5][0] ;
 wire \RAM[5][1] ;
 wire \RAM[5][2] ;
 wire \RAM[5][3] ;
 wire \RAM[5][4] ;
 wire \RAM[5][5] ;
 wire \RAM[61][0] ;
 wire \RAM[61][1] ;
 wire \RAM[61][2] ;
 wire \RAM[61][3] ;
 wire \RAM[61][4] ;
 wire \RAM[61][5] ;
 wire \RAM[62][0] ;
 wire \RAM[62][1] ;
 wire \RAM[62][2] ;
 wire \RAM[62][3] ;
 wire \RAM[62][4] ;
 wire \RAM[62][5] ;
 wire \RAM[6][0] ;
 wire \RAM[6][1] ;
 wire \RAM[6][2] ;
 wire \RAM[6][3] ;
 wire \RAM[6][4] ;
 wire \RAM[6][5] ;
 wire \RAM[7][0] ;
 wire \RAM[7][1] ;
 wire \RAM[7][2] ;
 wire \RAM[7][3] ;
 wire \RAM[7][4] ;
 wire \RAM[7][5] ;
 wire \RAM[8][0] ;
 wire \RAM[8][1] ;
 wire \RAM[8][2] ;
 wire \RAM[8][3] ;
 wire \RAM[8][4] ;
 wire \RAM[8][5] ;
 wire \RAM[9][0] ;
 wire \RAM[9][1] ;
 wire \RAM[9][2] ;
 wire \RAM[9][3] ;
 wire \RAM[9][4] ;
 wire \RAM[9][5] ;
 wire ROM_DO;
 wire \ROM_addr_buff[0] ;
 wire \ROM_addr_buff[10] ;
 wire \ROM_addr_buff[11] ;
 wire \ROM_addr_buff[1] ;
 wire \ROM_addr_buff[2] ;
 wire \ROM_addr_buff[3] ;
 wire \ROM_addr_buff[4] ;
 wire \ROM_addr_buff[5] ;
 wire \ROM_addr_buff[6] ;
 wire \ROM_addr_buff[7] ;
 wire \ROM_addr_buff[8] ;
 wire \ROM_addr_buff[9] ;
 wire \ROM_dest[0] ;
 wire \ROM_dest[1] ;
 wire \ROM_dest[2] ;
 wire \ROM_spi_cycle[0] ;
 wire \ROM_spi_cycle[1] ;
 wire \ROM_spi_cycle[2] ;
 wire \ROM_spi_cycle[3] ;
 wire \ROM_spi_cycle[4] ;
 wire \ROM_spi_dat_out[0] ;
 wire \ROM_spi_dat_out[1] ;
 wire \ROM_spi_dat_out[2] ;
 wire \ROM_spi_dat_out[3] ;
 wire \ROM_spi_dat_out[4] ;
 wire \ROM_spi_dat_out[5] ;
 wire \ROM_spi_dat_out[6] ;
 wire \ROM_spi_dat_out[7] ;
 wire SCLK_ROM;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire carry;
 wire compat;
 wire \imm_buff[0] ;
 wire \imm_buff[1] ;
 wire \imm_buff[2] ;
 wire \imm_buff[3] ;
 wire \imm_buff[4] ;
 wire \imm_buff[5] ;
 wire in_irupt;
 wire \insin[0] ;
 wire \insin[1] ;
 wire \insin[2] ;
 wire \insin[3] ;
 wire \insin[4] ;
 wire \insin[5] ;
 wire \instr_cycle[0] ;
 wire \instr_cycle[1] ;
 wire \instr_cycle[2] ;
 wire \last_A[0] ;
 wire \last_A[1] ;
 wire \last_A[2] ;
 wire \last_A[3] ;
 wire \last_A[4] ;
 wire \last_A[5] ;
 wire \last_B[0] ;
 wire \last_B[1] ;
 wire \last_B[2] ;
 wire \last_B[3] ;
 wire \last_B[4] ;
 wire \last_B[5] ;
 wire \last_MAR[0] ;
 wire \last_MAR[1] ;
 wire \last_MAR[2] ;
 wire \last_MAR[3] ;
 wire \last_MAR[4] ;
 wire \last_MAR[5] ;
 wire \last_PC[0] ;
 wire \last_PC[10] ;
 wire \last_PC[11] ;
 wire \last_PC[1] ;
 wire \last_PC[2] ;
 wire \last_PC[3] ;
 wire \last_PC[4] ;
 wire \last_PC[5] ;
 wire \last_PC[6] ;
 wire \last_PC[7] ;
 wire \last_PC[8] ;
 wire \last_PC[9] ;
 wire \last_P[0] ;
 wire \last_P[1] ;
 wire \last_P[2] ;
 wire \last_P[3] ;
 wire \last_P[4] ;
 wire \last_P[5] ;
 wire \last_addr[0] ;
 wire \last_addr[10] ;
 wire \last_addr[11] ;
 wire \last_addr[1] ;
 wire \last_addr[2] ;
 wire \last_addr[3] ;
 wire \last_addr[4] ;
 wire \last_addr[5] ;
 wire \last_addr[6] ;
 wire \last_addr[7] ;
 wire \last_addr[8] ;
 wire \last_addr[9] ;
 wire \last_flags[0] ;
 wire \last_flags[1] ;
 wire last_inter;
 wire \mem_cycle[0] ;
 wire \mem_cycle[1] ;
 wire \mem_cycle[2] ;
 wire needs_irupt;
 wire spi_clkdiv;
 wire net164;
 wire clknet_leaf_0_clk;
 wire net165;
 wire zero;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;

 sky130_as_sc_hs__inv_2 _2514_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\ROM_spi_cycle[1] ),
    .Y(_0526_));
 sky130_as_sc_hs__nor2_2 _2515_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\ROM_spi_cycle[3] ),
    .B(\ROM_spi_cycle[2] ),
    .Y(_0527_));
 sky130_as_sc_hs__and2_2 _2516_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0526_),
    .B(_0527_),
    .Y(_0528_));
 sky130_as_sc_hs__nor2_2 _2517_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\ROM_spi_cycle[4] ),
    .B(\ROM_spi_cycle[0] ),
    .Y(_0529_));
 sky130_as_sc_hs__nand2_4 _2518_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0528_),
    .B(_0529_),
    .Y(_0530_));
 sky130_as_sc_hs__or2_4 _2519_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net143),
    .B(\mem_cycle[1] ),
    .Y(_0531_));
 sky130_as_sc_hs__or2_2 _2520_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net144),
    .B(_0531_),
    .Y(_0532_));
 sky130_as_sc_hs__nor2_4 _2521_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0530_),
    .B(_0532_),
    .Y(_0533_));
 sky130_as_sc_hs__nor2_2 _2522_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net138),
    .B(net136),
    .Y(_0534_));
 sky130_as_sc_hs__inv_2 _2523_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net49),
    .Y(_0535_));
 sky130_as_sc_hs__mux2_2 _2524_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net93),
    .B(\RAM[22][2] ),
    .A(\RAM[20][2] ),
    .Y(_0536_));
 sky130_as_sc_hs__mux2_2 _2525_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net93),
    .B(\RAM[23][2] ),
    .A(\RAM[21][2] ),
    .Y(_0537_));
 sky130_as_sc_hs__mux2_2 _2526_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net119),
    .B(_0537_),
    .A(_0536_),
    .Y(_0538_));
 sky130_as_sc_hs__mux2_2 _2527_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net65),
    .B(\RAM[18][2] ),
    .A(\RAM[16][2] ),
    .Y(_0539_));
 sky130_as_sc_hs__mux2_2 _2528_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net65),
    .B(\RAM[19][2] ),
    .A(\RAM[17][2] ),
    .Y(_0540_));
 sky130_as_sc_hs__mux2_2 _2529_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net104),
    .B(_0540_),
    .A(_0539_),
    .Y(_0541_));
 sky130_as_sc_hs__inv_4 _2530_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net62),
    .Y(_0542_));
 sky130_as_sc_hs__mux2_2 _2531_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0542_),
    .B(_0541_),
    .A(_0538_),
    .Y(_0543_));
 sky130_as_sc_hs__mux2_2 _2532_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net92),
    .B(\RAM[30][2] ),
    .A(\RAM[28][2] ),
    .Y(_0544_));
 sky130_as_sc_hs__mux2_2 _2533_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net92),
    .B(\RAM[31][2] ),
    .A(\RAM[29][2] ),
    .Y(_0545_));
 sky130_as_sc_hs__mux2_2 _2534_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net119),
    .B(_0545_),
    .A(_0544_),
    .Y(_0546_));
 sky130_as_sc_hs__mux2_2 _2535_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net96),
    .B(\RAM[26][2] ),
    .A(\RAM[24][2] ),
    .Y(_0547_));
 sky130_as_sc_hs__mux2_2 _2536_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net97),
    .B(\RAM[27][2] ),
    .A(\RAM[25][2] ),
    .Y(_0548_));
 sky130_as_sc_hs__mux2_2 _2537_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net120),
    .B(_0548_),
    .A(_0547_),
    .Y(_0549_));
 sky130_as_sc_hs__mux2_2 _2538_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0542_),
    .B(_0549_),
    .A(_0546_),
    .Y(_0550_));
 sky130_as_sc_hs__mux2_2 _2539_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net54),
    .B(_0550_),
    .A(_0543_),
    .Y(_0551_));
 sky130_as_sc_hs__inv_2 _2540_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net54),
    .Y(_0552_));
 sky130_as_sc_hs__nor2_2 _2541_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0552_),
    .B(net141),
    .Y(_0553_));
 sky130_as_sc_hs__mux2_2 _2542_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net98),
    .B(\RAM[14][2] ),
    .A(\RAM[12][2] ),
    .Y(_0554_));
 sky130_as_sc_hs__mux2_2 _2543_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net98),
    .B(\RAM[15][2] ),
    .A(\RAM[13][2] ),
    .Y(_0555_));
 sky130_as_sc_hs__mux2_2 _2544_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net121),
    .B(_0555_),
    .A(_0554_),
    .Y(_0556_));
 sky130_as_sc_hs__mux2_2 _2545_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net98),
    .B(\RAM[10][2] ),
    .A(\RAM[8][2] ),
    .Y(_0557_));
 sky130_as_sc_hs__mux2_2 _2546_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net98),
    .B(\RAM[11][2] ),
    .A(\RAM[9][2] ),
    .Y(_0558_));
 sky130_as_sc_hs__mux2_2 _2547_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net120),
    .B(_0558_),
    .A(_0557_),
    .Y(_0559_));
 sky130_as_sc_hs__buff_6 _2548_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0542_),
    .Y(_0560_));
 sky130_as_sc_hs__mux2_2 _2549_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0560_),
    .B(_0559_),
    .A(_0556_),
    .Y(_0561_));
 sky130_as_sc_hs__nor2_2 _2550_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net54),
    .B(net141),
    .Y(_0562_));
 sky130_as_sc_hs__or2_2 _2551_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net57),
    .B(net68),
    .Y(_0563_));
 sky130_as_sc_hs__mux2_2 _2552_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net105),
    .B(\RAM[1][2] ),
    .A(\RAM[0][2] ),
    .Y(_0564_));
 sky130_as_sc_hs__nand2b_2 _2553_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(net73),
    .Y(_0565_),
    .A(net57));
 sky130_as_sc_hs__mux2_2 _2554_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net105),
    .B(\RAM[3][2] ),
    .A(\RAM[2][2] ),
    .Y(_0566_));
 sky130_as_sc_hs__oa22_2 _2555_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0563_),
    .B(_0564_),
    .C(_0565_),
    .D(_0566_),
    .Y(_0567_));
 sky130_as_sc_hs__nand2_2 _2556_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net58),
    .B(net84),
    .Y(_0568_));
 sky130_as_sc_hs__mux2_2 _2557_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net109),
    .B(\RAM[7][2] ),
    .A(\RAM[6][2] ),
    .Y(_0569_));
 sky130_as_sc_hs__mux2_2 _2558_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net109),
    .B(\RAM[5][2] ),
    .A(\RAM[4][2] ),
    .Y(_0570_));
 sky130_as_sc_hs__nand2b_2 _2559_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(net58),
    .Y(_0571_),
    .A(net84));
 sky130_as_sc_hs__oa22_2 _2560_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0568_),
    .B(_0569_),
    .C(_0570_),
    .D(_0571_),
    .Y(_0572_));
 sky130_as_sc_hs__nor2_2 _2561_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0535_),
    .B(net141),
    .Y(_0573_));
 sky130_as_sc_hs__ao31_2 _2562_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0562_),
    .B(_0567_),
    .C(_0572_),
    .D(_0573_),
    .Y(_0574_));
 sky130_as_sc_hs__ao21_2 _2563_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0553_),
    .B(_0561_),
    .C(_0574_),
    .Y(_0575_));
 sky130_as_sc_hs__oa21_2 _2564_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0535_),
    .B(_0551_),
    .C(_0575_),
    .Y(_0576_));
 sky130_as_sc_hs__or2_2 _2565_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net42),
    .B(net35),
    .Y(_0577_));
 sky130_as_sc_hs__nor3_2 _2566_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net39),
    .B(net47),
    .C(net29),
    .Y(_0578_));
 sky130_as_sc_hs__nor2b_2 _2567_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0577_),
    .Y(_0579_),
    .B(_0578_));
 sky130_as_sc_hs__nand4_2 _2568_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net39),
    .B(net47),
    .C(net40),
    .Y(_0580_),
    .D(net35));
 sky130_as_sc_hs__nand2_2 _2569_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net34),
    .B(net29),
    .Y(_0581_));
 sky130_as_sc_hs__nor2_2 _2570_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0580_),
    .B(_0581_),
    .Y(_0582_));
 sky130_as_sc_hs__nand2b_2 _2571_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(net40),
    .Y(_0583_),
    .A(net47));
 sky130_as_sc_hs__nand2_2 _2572_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net39),
    .B(net35),
    .Y(_0584_));
 sky130_as_sc_hs__aoi211_2 _2573_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_0583_),
    .C(_0584_),
    .D(net29),
    .Y(_0585_),
    .A(net31));
 sky130_as_sc_hs__aoi211_2 _2574_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_0579_),
    .C(_0582_),
    .D(_0585_),
    .Y(_0586_),
    .A(net31));
 sky130_as_sc_hs__buff_4 _2575_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net23),
    .Y(_0587_));
 sky130_as_sc_hs__inv_2 _2576_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net140),
    .Y(_0588_));
 sky130_as_sc_hs__or2_2 _2577_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net52),
    .B(net49),
    .Y(_0589_));
 sky130_as_sc_hs__nor2_2 _2578_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0588_),
    .B(_0589_),
    .Y(_0590_));
 sky130_as_sc_hs__mux2_2 _2579_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net68),
    .B(\RAM[38][2] ),
    .A(\RAM[36][2] ),
    .Y(_0591_));
 sky130_as_sc_hs__mux2_2 _2580_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net68),
    .B(\RAM[39][2] ),
    .A(\RAM[37][2] ),
    .Y(_0592_));
 sky130_as_sc_hs__mux2_2 _2581_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net107),
    .B(_0592_),
    .A(_0591_),
    .Y(_0593_));
 sky130_as_sc_hs__mux2_2 _2582_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net64),
    .B(\RAM[34][2] ),
    .A(\RAM[32][2] ),
    .Y(_0594_));
 sky130_as_sc_hs__mux2_2 _2583_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net64),
    .B(\RAM[35][2] ),
    .A(\RAM[33][2] ),
    .Y(_0595_));
 sky130_as_sc_hs__mux2_2 _2584_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net104),
    .B(_0595_),
    .A(_0594_),
    .Y(_0596_));
 sky130_as_sc_hs__buff_6 _2585_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0542_),
    .Y(_0597_));
 sky130_as_sc_hs__mux2_2 _2586_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0597_),
    .B(_0596_),
    .A(_0593_),
    .Y(_0598_));
 sky130_as_sc_hs__mux2_2 _2587_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net86),
    .B(\RAM[62][2] ),
    .A(uo_out[2]),
    .Y(_0599_));
 sky130_as_sc_hs__mux2_2 _2588_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net81),
    .B(uio_out[2]),
    .A(\RAM[61][2] ),
    .Y(_0600_));
 sky130_as_sc_hs__mux2_2 _2589_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net116),
    .B(_0600_),
    .A(_0599_),
    .Y(_0601_));
 sky130_as_sc_hs__mux2_2 _2590_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net87),
    .B(\RAM[58][2] ),
    .A(\RAM[56][2] ),
    .Y(_0602_));
 sky130_as_sc_hs__mux2_2 _2591_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net80),
    .B(uio_oe[2]),
    .A(\RAM[57][2] ),
    .Y(_0603_));
 sky130_as_sc_hs__mux2_2 _2592_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net116),
    .B(_0603_),
    .A(_0602_),
    .Y(_0604_));
 sky130_as_sc_hs__mux2_2 _2593_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0597_),
    .B(_0604_),
    .A(_0601_),
    .Y(_0605_));
 sky130_as_sc_hs__nand2_2 _2594_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net52),
    .B(net49),
    .Y(_0606_));
 sky130_as_sc_hs__nor2_4 _2595_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0588_),
    .B(_0606_),
    .Y(_0607_));
 sky130_as_sc_hs__aoi22_2 _2596_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0590_),
    .B(_0598_),
    .C(_0605_),
    .D(_0607_),
    .Y(_0608_));
 sky130_as_sc_hs__nand2b_2 _2597_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(net49),
    .Y(_0609_),
    .A(net52));
 sky130_as_sc_hs__nor2_2 _2598_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0588_),
    .B(_0609_),
    .Y(_0610_));
 sky130_as_sc_hs__mux2_2 _2599_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net77),
    .B(\RAM[54][2] ),
    .A(\RAM[52][2] ),
    .Y(_0611_));
 sky130_as_sc_hs__mux2_2 _2600_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net77),
    .B(\RAM[55][2] ),
    .A(\RAM[53][2] ),
    .Y(_0612_));
 sky130_as_sc_hs__mux2_2 _2601_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net112),
    .B(_0612_),
    .A(_0611_),
    .Y(_0613_));
 sky130_as_sc_hs__mux2_2 _2602_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net77),
    .B(\RAM[50][2] ),
    .A(\RAM[48][2] ),
    .Y(_0614_));
 sky130_as_sc_hs__mux2_2 _2603_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net83),
    .B(\RAM[51][2] ),
    .A(\RAM[49][2] ),
    .Y(_0615_));
 sky130_as_sc_hs__mux2_2 _2604_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net112),
    .B(_0615_),
    .A(_0614_),
    .Y(_0616_));
 sky130_as_sc_hs__mux2_2 _2605_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0597_),
    .B(_0616_),
    .A(_0613_),
    .Y(_0617_));
 sky130_as_sc_hs__nand2_2 _2606_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0610_),
    .B(_0617_),
    .Y(_0618_));
 sky130_as_sc_hs__inv_2 _2607_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net114),
    .Y(_0619_));
 sky130_as_sc_hs__buff_8 _2608_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0619_),
    .Y(_0620_));
 sky130_as_sc_hs__mux2_2 _2609_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net83),
    .B(\RAM[43][2] ),
    .A(\RAM[41][2] ),
    .Y(_0621_));
 sky130_as_sc_hs__mux2_2 _2610_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net80),
    .B(\RAM[47][2] ),
    .A(\RAM[45][2] ),
    .Y(_0622_));
 sky130_as_sc_hs__mux2_2 _2611_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net60),
    .B(_0622_),
    .A(_0621_),
    .Y(_0623_));
 sky130_as_sc_hs__nor2_2 _2612_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0620_),
    .B(_0623_),
    .Y(_0624_));
 sky130_as_sc_hs__or2_2 _2613_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net114),
    .B(net58),
    .Y(_0625_));
 sky130_as_sc_hs__mux2_2 _2614_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net75),
    .B(\RAM[42][2] ),
    .A(\RAM[40][2] ),
    .Y(_0626_));
 sky130_as_sc_hs__nand2b_2 _2615_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(net58),
    .Y(_0627_),
    .A(net115));
 sky130_as_sc_hs__mux2_2 _2616_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net78),
    .B(\RAM[46][2] ),
    .A(\RAM[44][2] ),
    .Y(_0628_));
 sky130_as_sc_hs__or2_2 _2617_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0627_),
    .B(_0628_),
    .Y(_0629_));
 sky130_as_sc_hs__nand2b_2 _2618_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(net52),
    .Y(_0630_),
    .A(net50));
 sky130_as_sc_hs__clkbuff_4 _2619_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0630_),
    .Y(_0631_));
 sky130_as_sc_hs__nor2_2 _2620_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0588_),
    .B(_0631_),
    .Y(_0632_));
 sky130_as_sc_hs__iao211_2 _2621_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0625_),
    .B(_0626_),
    .C(_0629_),
    .D(_0632_),
    .Y(_0633_));
 sky130_as_sc_hs__xnor2_2 _2622_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net114),
    .Y(_0634_),
    .B(net84));
 sky130_as_sc_hs__nand3_2 _2623_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net58),
    .B(_0607_),
    .C(_0634_),
    .Y(_0635_));
 sky130_as_sc_hs__oa21_2 _2624_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0624_),
    .B(_0633_),
    .C(_0635_),
    .Y(_0636_));
 sky130_as_sc_hs__nand4_2 _2625_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0587_),
    .B(_0608_),
    .C(_0618_),
    .Y(_0637_),
    .D(_0636_));
 sky130_as_sc_hs__nand3_2 _2626_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net53),
    .B(net50),
    .C(net140),
    .Y(_0638_));
 sky130_as_sc_hs__nand3_2 _2627_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net115),
    .B(net59),
    .C(net101),
    .Y(_0639_));
 sky130_as_sc_hs__or2_2 _2628_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_as_sc_hs__and2_2 _2629_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net52),
    .B(net49),
    .Y(_0641_));
 sky130_as_sc_hs__nor2b_2 _2630_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net101),
    .Y(_0642_),
    .B(net58));
 sky130_as_sc_hs__nand4_2 _2631_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net140),
    .B(_0620_),
    .C(_0641_),
    .Y(_0643_),
    .D(_0642_));
 sky130_as_sc_hs__oa22_2 _2632_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net12),
    .B(_0640_),
    .C(_0643_),
    .D(net4),
    .Y(_0644_));
 sky130_as_sc_hs__mux2_2 _2633_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0587_),
    .B(_0644_),
    .A(\imm_buff[2] ),
    .Y(_0645_));
 sky130_as_sc_hs__oa21_2 _2634_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0576_),
    .B(_0637_),
    .C(_0645_),
    .Y(_0646_));
 sky130_as_sc_hs__buff_4 _2635_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0646_),
    .Y(_0647_));
 sky130_as_sc_hs__inv_2 _2636_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net40),
    .Y(_0648_));
 sky130_as_sc_hs__nand2_4 _2637_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net37),
    .B(net45),
    .Y(_0649_));
 sky130_as_sc_hs__nor2_2 _2638_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0648_),
    .B(_0649_),
    .Y(_0650_));
 sky130_as_sc_hs__buff_4 _2639_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0650_),
    .Y(_0651_));
 sky130_as_sc_hs__nor2_2 _2640_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net33),
    .B(net36),
    .Y(_0652_));
 sky130_as_sc_hs__nand3_2 _2641_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\instr_cycle[1] ),
    .B(_0651_),
    .C(_0652_),
    .Y(_0653_));
 sky130_as_sc_hs__mux2_2 _2642_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0653_),
    .B(net61),
    .A(_0647_),
    .Y(_0654_));
 sky130_as_sc_hs__inv_2 _2643_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net136),
    .Y(_0655_));
 sky130_as_sc_hs__buff_4 _2644_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0655_),
    .Y(_0656_));
 sky130_as_sc_hs__nor2_2 _2645_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net138),
    .B(_0656_),
    .Y(_0657_));
 sky130_as_sc_hs__or2_2 _2646_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net38),
    .B(net35),
    .Y(_0658_));
 sky130_as_sc_hs__nor3_2 _2647_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0583_),
    .B(_0581_),
    .C(_0658_),
    .Y(_0659_));
 sky130_as_sc_hs__clkbuff_4 _2648_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0659_),
    .Y(_0660_));
 sky130_as_sc_hs__mux2_2 _2649_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0660_),
    .B(\last_MAR[2] ),
    .A(net61),
    .Y(_0661_));
 sky130_as_sc_hs__ao22_2 _2650_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0534_),
    .C(_0657_),
    .B(_0654_),
    .D(_0661_),
    .Y(_0662_));
 sky130_as_sc_hs__inv_2 _2651_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net139),
    .Y(_0663_));
 sky130_as_sc_hs__nand2_2 _2652_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0663_),
    .B(_0533_),
    .Y(_0664_));
 sky130_as_sc_hs__clkbuff_4 _2653_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0664_),
    .Y(_0665_));
 sky130_as_sc_hs__ao22_2 _2654_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0533_),
    .C(_0665_),
    .B(_0662_),
    .D(net63),
    .Y(_0666_));
 sky130_as_sc_hs__inv_2 _2655_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\ROM_dest[2] ),
    .Y(_0667_));
 sky130_as_sc_hs__and2_2 _2656_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0528_),
    .B(_0529_),
    .Y(_0668_));
 sky130_as_sc_hs__nand4_2 _2657_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net143),
    .B(\mem_cycle[1] ),
    .C(net144),
    .Y(_0669_),
    .D(_0668_));
 sky130_as_sc_hs__or2_2 _2658_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_dest[0] ),
    .B(_0669_),
    .Y(_0670_));
 sky130_as_sc_hs__or2_2 _2659_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0667_),
    .B(_0670_),
    .Y(_0671_));
 sky130_as_sc_hs__clkbuff_4 _2660_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0671_),
    .Y(_0672_));
 sky130_as_sc_hs__mux2_2 _2661_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0672_),
    .B(_0666_),
    .A(\ROM_spi_dat_out[2] ),
    .Y(_0673_));
 sky130_as_sc_hs__and2_2 _2662_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net149),
    .B(_0673_),
    .Y(_0674_));
 sky130_as_sc_hs__buff_2 _2663_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0674_),
    .Y(_0002_));
 sky130_as_sc_hs__buff_2 _2664_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0534_),
    .Y(_0675_));
 sky130_as_sc_hs__mux2_2 _2665_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net69),
    .B(\RAM[18][3] ),
    .A(\RAM[16][3] ),
    .Y(_0676_));
 sky130_as_sc_hs__mux2_2 _2666_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net67),
    .B(\RAM[19][3] ),
    .A(\RAM[17][3] ),
    .Y(_0677_));
 sky130_as_sc_hs__mux2_2 _2667_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net106),
    .B(_0677_),
    .A(_0676_),
    .Y(_0678_));
 sky130_as_sc_hs__nor2_2 _2668_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0535_),
    .B(net57),
    .Y(_0679_));
 sky130_as_sc_hs__mux2_2 _2669_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net70),
    .B(\RAM[2][3] ),
    .A(\RAM[0][3] ),
    .Y(_0680_));
 sky130_as_sc_hs__mux2_2 _2670_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net66),
    .B(\RAM[3][3] ),
    .A(\RAM[1][3] ),
    .Y(_0681_));
 sky130_as_sc_hs__mux2_2 _2671_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net109),
    .B(_0681_),
    .A(_0680_),
    .Y(_0682_));
 sky130_as_sc_hs__nor2_2 _2672_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net51),
    .B(net56),
    .Y(_0683_));
 sky130_as_sc_hs__nor2_2 _2673_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net51),
    .B(_0542_),
    .Y(_0684_));
 sky130_as_sc_hs__mux2_2 _2674_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net72),
    .B(\RAM[6][3] ),
    .A(\RAM[4][3] ),
    .Y(_0685_));
 sky130_as_sc_hs__mux2_2 _2675_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net90),
    .B(\RAM[7][3] ),
    .A(\RAM[5][3] ),
    .Y(_0686_));
 sky130_as_sc_hs__mux2_2 _2676_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net109),
    .B(_0686_),
    .A(_0685_),
    .Y(_0687_));
 sky130_as_sc_hs__ao22_2 _2677_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0682_),
    .C(_0684_),
    .B(_0683_),
    .D(_0687_),
    .Y(_0688_));
 sky130_as_sc_hs__ao21_2 _2678_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0678_),
    .B(_0679_),
    .C(_0688_),
    .Y(_0689_));
 sky130_as_sc_hs__mux2_2 _2679_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net93),
    .B(\RAM[22][3] ),
    .A(\RAM[20][3] ),
    .Y(_0690_));
 sky130_as_sc_hs__mux2_2 _2680_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net93),
    .B(\RAM[23][3] ),
    .A(\RAM[21][3] ),
    .Y(_0691_));
 sky130_as_sc_hs__mux2_2 _2681_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net119),
    .B(_0691_),
    .A(_0690_),
    .Y(_0692_));
 sky130_as_sc_hs__ao31_2 _2682_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net51),
    .B(net62),
    .C(_0692_),
    .D(net54),
    .Y(_0693_));
 sky130_as_sc_hs__and2_2 _2683_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net122),
    .B(net59),
    .Y(_0694_));
 sky130_as_sc_hs__buff_4 _2684_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0694_),
    .Y(_0695_));
 sky130_as_sc_hs__mux2_2 _2685_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net91),
    .B(\RAM[31][3] ),
    .A(\RAM[29][3] ),
    .Y(_0696_));
 sky130_as_sc_hs__mux2_2 _2686_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net90),
    .B(\RAM[27][3] ),
    .A(\RAM[25][3] ),
    .Y(_0697_));
 sky130_as_sc_hs__nor2b_2 _2687_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net61),
    .Y(_0698_),
    .B(net122));
 sky130_as_sc_hs__ao22_2 _2688_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0695_),
    .C(_0697_),
    .B(_0696_),
    .D(net26),
    .Y(_0699_));
 sky130_as_sc_hs__nor2b_2 _2689_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net122),
    .Y(_0700_),
    .B(net61));
 sky130_as_sc_hs__mux2_2 _2690_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net90),
    .B(\RAM[30][3] ),
    .A(\RAM[28][3] ),
    .Y(_0701_));
 sky130_as_sc_hs__mux2_2 _2691_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net91),
    .B(\RAM[26][3] ),
    .A(\RAM[24][3] ),
    .Y(_0702_));
 sky130_as_sc_hs__nor2_4 _2692_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net122),
    .B(net61),
    .Y(_0703_));
 sky130_as_sc_hs__ao22_2 _2693_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net25),
    .C(_0702_),
    .B(_0701_),
    .D(_0703_),
    .Y(_0704_));
 sky130_as_sc_hs__nor2_2 _2694_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0699_),
    .B(_0704_),
    .Y(_0705_));
 sky130_as_sc_hs__mux2_2 _2695_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net94),
    .B(\RAM[14][3] ),
    .A(\RAM[12][3] ),
    .Y(_0706_));
 sky130_as_sc_hs__mux2_2 _2696_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net94),
    .B(\RAM[15][3] ),
    .A(\RAM[13][3] ),
    .Y(_0707_));
 sky130_as_sc_hs__ao22_2 _2697_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net25),
    .C(_0707_),
    .B(_0706_),
    .D(_0695_),
    .Y(_0708_));
 sky130_as_sc_hs__mux2_2 _2698_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net91),
    .B(\RAM[10][3] ),
    .A(\RAM[8][3] ),
    .Y(_0709_));
 sky130_as_sc_hs__mux2_2 _2699_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net94),
    .B(\RAM[11][3] ),
    .A(\RAM[9][3] ),
    .Y(_0710_));
 sky130_as_sc_hs__ao22_2 _2700_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0703_),
    .C(net26),
    .B(_0709_),
    .D(_0710_),
    .Y(_0711_));
 sky130_as_sc_hs__nor3_2 _2701_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0631_),
    .B(_0708_),
    .C(_0711_),
    .Y(_0712_));
 sky130_as_sc_hs__aoi211_2 _2702_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_0705_),
    .C(_0712_),
    .D(net141),
    .Y(_0713_),
    .A(_0641_));
 sky130_as_sc_hs__oai21_2 _2703_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0689_),
    .B(_0693_),
    .C(_0713_),
    .Y(_0714_));
 sky130_as_sc_hs__mux2_2 _2704_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net80),
    .B(\RAM[43][3] ),
    .A(\RAM[41][3] ),
    .Y(_0715_));
 sky130_as_sc_hs__mux2_2 _2705_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net80),
    .B(\RAM[47][3] ),
    .A(\RAM[45][3] ),
    .Y(_0716_));
 sky130_as_sc_hs__mux2_2 _2706_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net60),
    .B(_0716_),
    .A(_0715_),
    .Y(_0717_));
 sky130_as_sc_hs__mux2_2 _2707_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net80),
    .B(\RAM[42][3] ),
    .A(\RAM[40][3] ),
    .Y(_0718_));
 sky130_as_sc_hs__mux2_2 _2708_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net78),
    .B(\RAM[46][3] ),
    .A(\RAM[44][3] ),
    .Y(_0719_));
 sky130_as_sc_hs__mux2_2 _2709_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net60),
    .B(_0719_),
    .A(_0718_),
    .Y(_0720_));
 sky130_as_sc_hs__mux2_2 _2710_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0620_),
    .B(_0720_),
    .A(_0717_),
    .Y(_0721_));
 sky130_as_sc_hs__mux2_2 _2711_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net68),
    .B(\RAM[38][3] ),
    .A(\RAM[36][3] ),
    .Y(_0722_));
 sky130_as_sc_hs__mux2_2 _2712_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net68),
    .B(\RAM[39][3] ),
    .A(\RAM[37][3] ),
    .Y(_0723_));
 sky130_as_sc_hs__mux2_2 _2713_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net106),
    .B(_0723_),
    .A(_0722_),
    .Y(_0724_));
 sky130_as_sc_hs__mux2_2 _2714_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net64),
    .B(\RAM[34][3] ),
    .A(\RAM[32][3] ),
    .Y(_0725_));
 sky130_as_sc_hs__mux2_2 _2715_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net64),
    .B(\RAM[35][3] ),
    .A(\RAM[33][3] ),
    .Y(_0726_));
 sky130_as_sc_hs__mux2_2 _2716_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net104),
    .B(_0726_),
    .A(_0725_),
    .Y(_0727_));
 sky130_as_sc_hs__mux2_2 _2717_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0560_),
    .B(_0727_),
    .A(_0724_),
    .Y(_0728_));
 sky130_as_sc_hs__oa22_2 _2718_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0631_),
    .B(_0721_),
    .C(_0728_),
    .D(_0589_),
    .Y(_0729_));
 sky130_as_sc_hs__mux2_2 _2719_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net86),
    .B(\RAM[62][3] ),
    .A(uo_out[3]),
    .Y(_0730_));
 sky130_as_sc_hs__aoi21_2 _2720_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0700_),
    .B(_0730_),
    .C(_0606_),
    .Y(_0731_));
 sky130_as_sc_hs__mux2_2 _2721_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net81),
    .B(uio_out[3]),
    .A(\RAM[61][3] ),
    .Y(_0732_));
 sky130_as_sc_hs__mux2_2 _2722_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net86),
    .B(uio_oe[3]),
    .A(\RAM[57][3] ),
    .Y(_0733_));
 sky130_as_sc_hs__mux2_2 _2723_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net101),
    .B(\RAM[58][3] ),
    .A(\RAM[56][3] ),
    .Y(_0734_));
 sky130_as_sc_hs__ao22_2 _2724_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0698_),
    .C(_0734_),
    .B(_0733_),
    .D(_0703_),
    .Y(_0735_));
 sky130_as_sc_hs__aoi21_2 _2725_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0695_),
    .B(_0732_),
    .C(_0735_),
    .Y(_0736_));
 sky130_as_sc_hs__ao31_2 _2726_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0619_),
    .B(_0641_),
    .C(_0642_),
    .D(_0588_),
    .Y(_0737_));
 sky130_as_sc_hs__mux2_2 _2727_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net106),
    .B(\RAM[49][3] ),
    .A(\RAM[48][3] ),
    .Y(_0738_));
 sky130_as_sc_hs__mux2_2 _2728_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net107),
    .B(\RAM[51][3] ),
    .A(\RAM[50][3] ),
    .Y(_0739_));
 sky130_as_sc_hs__oa22_2 _2729_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0563_),
    .B(_0738_),
    .C(_0739_),
    .D(_0565_),
    .Y(_0740_));
 sky130_as_sc_hs__mux2_2 _2730_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net113),
    .B(\RAM[53][3] ),
    .A(\RAM[52][3] ),
    .Y(_0741_));
 sky130_as_sc_hs__mux2_2 _2731_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net114),
    .B(\RAM[55][3] ),
    .A(\RAM[54][3] ),
    .Y(_0742_));
 sky130_as_sc_hs__oa22_2 _2732_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0571_),
    .B(_0741_),
    .C(_0742_),
    .D(_0568_),
    .Y(_0743_));
 sky130_as_sc_hs__aoi21_2 _2733_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0740_),
    .B(_0743_),
    .C(_0609_),
    .Y(_0744_));
 sky130_as_sc_hs__aoi211_2 _2734_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_0736_),
    .C(_0737_),
    .D(_0744_),
    .Y(_0745_),
    .A(_0731_));
 sky130_as_sc_hs__nor3_2 _2735_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net114),
    .B(_0638_),
    .C(_0571_),
    .Y(_0746_));
 sky130_as_sc_hs__nor2_2 _2736_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0638_),
    .B(_0639_),
    .Y(_0747_));
 sky130_as_sc_hs__ao21_2 _2737_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net5),
    .B(net24),
    .C(_0747_),
    .Y(_0748_));
 sky130_as_sc_hs__aoi21_2 _2738_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0729_),
    .B(_0745_),
    .C(_0748_),
    .Y(_0749_));
 sky130_as_sc_hs__inv_2 _2739_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net13),
    .Y(_0750_));
 sky130_as_sc_hs__nor2_2 _2740_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\imm_buff[3] ),
    .B(_0587_),
    .Y(_0751_));
 sky130_as_sc_hs__ao31_2 _2741_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0750_),
    .B(_0586_),
    .C(_0747_),
    .D(_0751_),
    .Y(_0752_));
 sky130_as_sc_hs__ao31_4 _2742_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0587_),
    .B(_0714_),
    .C(_0749_),
    .D(_0752_),
    .Y(_0753_));
 sky130_as_sc_hs__buff_8 _2743_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0753_),
    .Y(_0754_));
 sky130_as_sc_hs__nand2_2 _2744_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net53),
    .B(_0653_),
    .Y(_0755_));
 sky130_as_sc_hs__oai21_2 _2745_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0653_),
    .B(_0754_),
    .C(_0755_),
    .Y(_0756_));
 sky130_as_sc_hs__buff_4 _2746_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0660_),
    .Y(_0757_));
 sky130_as_sc_hs__mux2_2 _2747_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0757_),
    .B(\last_MAR[3] ),
    .A(net53),
    .Y(_0758_));
 sky130_as_sc_hs__buff_2 _2748_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0657_),
    .Y(_0759_));
 sky130_as_sc_hs__ao22_2 _2749_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0675_),
    .C(_0758_),
    .B(_0756_),
    .D(_0759_),
    .Y(_0760_));
 sky130_as_sc_hs__clkbuff_4 _2750_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0533_),
    .Y(_0761_));
 sky130_as_sc_hs__ao22_2 _2751_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net53),
    .C(_0760_),
    .B(_0665_),
    .D(_0761_),
    .Y(_0762_));
 sky130_as_sc_hs__mux2_2 _2752_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0672_),
    .B(_0762_),
    .A(\ROM_spi_dat_out[3] ),
    .Y(_0763_));
 sky130_as_sc_hs__and2_2 _2753_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net149),
    .B(_0763_),
    .Y(_0764_));
 sky130_as_sc_hs__buff_2 _2754_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0764_),
    .Y(_0003_));
 sky130_as_sc_hs__mux2_2 _2755_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net68),
    .B(\RAM[38][4] ),
    .A(\RAM[36][4] ),
    .Y(_0765_));
 sky130_as_sc_hs__mux2_2 _2756_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net67),
    .B(\RAM[39][4] ),
    .A(\RAM[37][4] ),
    .Y(_0766_));
 sky130_as_sc_hs__mux2_2 _2757_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net106),
    .B(_0766_),
    .A(_0765_),
    .Y(_0767_));
 sky130_as_sc_hs__mux2_2 _2758_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net66),
    .B(\RAM[34][4] ),
    .A(\RAM[32][4] ),
    .Y(_0768_));
 sky130_as_sc_hs__mux2_2 _2759_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net66),
    .B(\RAM[35][4] ),
    .A(\RAM[33][4] ),
    .Y(_0769_));
 sky130_as_sc_hs__mux2_2 _2760_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net105),
    .B(_0769_),
    .A(_0768_),
    .Y(_0770_));
 sky130_as_sc_hs__mux2_2 _2761_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0560_),
    .B(_0770_),
    .A(_0767_),
    .Y(_0771_));
 sky130_as_sc_hs__mux2_2 _2762_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net79),
    .B(\RAM[46][4] ),
    .A(\RAM[44][4] ),
    .Y(_0772_));
 sky130_as_sc_hs__mux2_2 _2763_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net79),
    .B(\RAM[47][4] ),
    .A(\RAM[45][4] ),
    .Y(_0773_));
 sky130_as_sc_hs__mux2_2 _2764_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net117),
    .B(_0773_),
    .A(_0772_),
    .Y(_0774_));
 sky130_as_sc_hs__mux2_2 _2765_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net78),
    .B(\RAM[42][4] ),
    .A(\RAM[40][4] ),
    .Y(_0775_));
 sky130_as_sc_hs__mux2_2 _2766_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net78),
    .B(\RAM[43][4] ),
    .A(\RAM[41][4] ),
    .Y(_0776_));
 sky130_as_sc_hs__mux2_2 _2767_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net113),
    .B(_0776_),
    .A(_0775_),
    .Y(_0777_));
 sky130_as_sc_hs__mux2_2 _2768_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0597_),
    .B(_0777_),
    .A(_0774_),
    .Y(_0778_));
 sky130_as_sc_hs__mux2_2 _2769_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net55),
    .B(_0778_),
    .A(_0771_),
    .Y(_0779_));
 sky130_as_sc_hs__and2_2 _2770_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net31),
    .B(_0583_),
    .Y(_0780_));
 sky130_as_sc_hs__or2_2 _2771_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net29),
    .B(_0584_),
    .Y(_0781_));
 sky130_as_sc_hs__or2_2 _2772_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0580_),
    .B(_0581_),
    .Y(_0782_));
 sky130_as_sc_hs__inv_2 _2773_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net35),
    .Y(_0783_));
 sky130_as_sc_hs__nand4_2 _2774_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net31),
    .B(_0648_),
    .C(_0783_),
    .Y(_0784_),
    .D(_0578_));
 sky130_as_sc_hs__iao211_2 _2775_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0780_),
    .B(_0781_),
    .C(_0782_),
    .D(_0784_),
    .Y(_0785_));
 sky130_as_sc_hs__ao21_2 _2776_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\imm_buff[4] ),
    .B(net22),
    .C(_0747_),
    .Y(_0786_));
 sky130_as_sc_hs__aoi31_2 _2777_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0535_),
    .B(net140),
    .C(_0779_),
    .D(_0786_),
    .Y(_0787_));
 sky130_as_sc_hs__nor2_2 _2778_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net51),
    .B(net141),
    .Y(_0788_));
 sky130_as_sc_hs__mux2_2 _2779_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net71),
    .B(\RAM[30][4] ),
    .A(\RAM[28][4] ),
    .Y(_0789_));
 sky130_as_sc_hs__mux2_2 _2780_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net71),
    .B(\RAM[31][4] ),
    .A(\RAM[29][4] ),
    .Y(_0790_));
 sky130_as_sc_hs__mux2_2 _2781_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net111),
    .B(_0790_),
    .A(_0789_),
    .Y(_0791_));
 sky130_as_sc_hs__mux2_2 _2782_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net96),
    .B(\RAM[26][4] ),
    .A(\RAM[24][4] ),
    .Y(_0792_));
 sky130_as_sc_hs__mux2_2 _2783_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net96),
    .B(\RAM[27][4] ),
    .A(\RAM[25][4] ),
    .Y(_0793_));
 sky130_as_sc_hs__mux2_2 _2784_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net120),
    .B(_0793_),
    .A(_0792_),
    .Y(_0794_));
 sky130_as_sc_hs__mux2_2 _2785_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0597_),
    .B(_0794_),
    .A(_0791_),
    .Y(_0795_));
 sky130_as_sc_hs__mux2_2 _2786_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net56),
    .B(\RAM[20][4] ),
    .A(\RAM[16][4] ),
    .Y(_0796_));
 sky130_as_sc_hs__mux2_2 _2787_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net56),
    .B(\RAM[21][4] ),
    .A(\RAM[17][4] ),
    .Y(_0797_));
 sky130_as_sc_hs__mux2_2 _2788_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net110),
    .B(_0797_),
    .A(_0796_),
    .Y(_0798_));
 sky130_as_sc_hs__mux2_2 _2789_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net56),
    .B(\RAM[22][4] ),
    .A(\RAM[18][4] ),
    .Y(_0799_));
 sky130_as_sc_hs__mux2_2 _2790_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net56),
    .B(\RAM[23][4] ),
    .A(\RAM[19][4] ),
    .Y(_0800_));
 sky130_as_sc_hs__mux2_2 _2791_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net110),
    .B(_0800_),
    .A(_0799_),
    .Y(_0801_));
 sky130_as_sc_hs__mux2_2 _2792_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net73),
    .B(_0801_),
    .A(_0798_),
    .Y(_0802_));
 sky130_as_sc_hs__ao22_2 _2793_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0553_),
    .C(_0802_),
    .B(_0795_),
    .D(_0562_),
    .Y(_0803_));
 sky130_as_sc_hs__mux2_2 _2794_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net100),
    .B(\RAM[11][4] ),
    .A(\RAM[9][4] ),
    .Y(_0804_));
 sky130_as_sc_hs__mux2_2 _2795_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net99),
    .B(\RAM[15][4] ),
    .A(\RAM[13][4] ),
    .Y(_0805_));
 sky130_as_sc_hs__mux2_2 _2796_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net62),
    .B(_0805_),
    .A(_0804_),
    .Y(_0806_));
 sky130_as_sc_hs__mux2_2 _2797_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net96),
    .B(\RAM[10][4] ),
    .A(\RAM[8][4] ),
    .Y(_0807_));
 sky130_as_sc_hs__mux2_2 _2798_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net99),
    .B(\RAM[14][4] ),
    .A(\RAM[12][4] ),
    .Y(_0808_));
 sky130_as_sc_hs__mux2_2 _2799_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net62),
    .B(_0808_),
    .A(_0807_),
    .Y(_0809_));
 sky130_as_sc_hs__mux2_2 _2800_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0620_),
    .B(_0809_),
    .A(_0806_),
    .Y(_0810_));
 sky130_as_sc_hs__mux2_2 _2801_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net72),
    .B(\RAM[6][4] ),
    .A(\RAM[4][4] ),
    .Y(_0811_));
 sky130_as_sc_hs__mux2_2 _2802_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net90),
    .B(\RAM[7][4] ),
    .A(\RAM[5][4] ),
    .Y(_0812_));
 sky130_as_sc_hs__mux2_2 _2803_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net111),
    .B(_0812_),
    .A(_0811_),
    .Y(_0813_));
 sky130_as_sc_hs__mux2_2 _2804_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net70),
    .B(\RAM[2][4] ),
    .A(\RAM[0][4] ),
    .Y(_0814_));
 sky130_as_sc_hs__mux2_2 _2805_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net66),
    .B(\RAM[3][4] ),
    .A(\RAM[1][4] ),
    .Y(_0815_));
 sky130_as_sc_hs__mux2_2 _2806_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net105),
    .B(_0815_),
    .A(_0814_),
    .Y(_0816_));
 sky130_as_sc_hs__mux2_2 _2807_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0560_),
    .B(_0816_),
    .A(_0813_),
    .Y(_0817_));
 sky130_as_sc_hs__mux2_2 _2808_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0552_),
    .B(_0817_),
    .A(_0810_),
    .Y(_0818_));
 sky130_as_sc_hs__oai22_2 _2809_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0788_),
    .B(_0803_),
    .C(_0818_),
    .D(net51),
    .Y(_0819_));
 sky130_as_sc_hs__mux2_2 _2810_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net86),
    .B(\RAM[62][4] ),
    .A(uo_out[4]),
    .Y(_0820_));
 sky130_as_sc_hs__mux2_2 _2811_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net80),
    .B(uio_out[4]),
    .A(\RAM[61][4] ),
    .Y(_0821_));
 sky130_as_sc_hs__mux2_2 _2812_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net113),
    .B(_0821_),
    .A(_0820_),
    .Y(_0822_));
 sky130_as_sc_hs__mux2_2 _2813_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net101),
    .B(\RAM[58][4] ),
    .A(\RAM[56][4] ),
    .Y(_0823_));
 sky130_as_sc_hs__mux2_2 _2814_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net80),
    .B(uio_oe[4]),
    .A(\RAM[57][4] ),
    .Y(_0824_));
 sky130_as_sc_hs__mux2_2 _2815_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net113),
    .B(_0824_),
    .A(_0823_),
    .Y(_0825_));
 sky130_as_sc_hs__mux2_2 _2816_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0560_),
    .B(_0825_),
    .A(_0822_),
    .Y(_0826_));
 sky130_as_sc_hs__mux2_2 _2817_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net75),
    .B(\RAM[54][4] ),
    .A(\RAM[52][4] ),
    .Y(_0827_));
 sky130_as_sc_hs__mux2_2 _2818_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net76),
    .B(\RAM[55][4] ),
    .A(\RAM[53][4] ),
    .Y(_0828_));
 sky130_as_sc_hs__mux2_2 _2819_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net112),
    .B(_0828_),
    .A(_0827_),
    .Y(_0829_));
 sky130_as_sc_hs__mux2_2 _2820_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net75),
    .B(\RAM[50][4] ),
    .A(\RAM[48][4] ),
    .Y(_0830_));
 sky130_as_sc_hs__mux2_2 _2821_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net75),
    .B(\RAM[51][4] ),
    .A(\RAM[49][4] ),
    .Y(_0831_));
 sky130_as_sc_hs__mux2_2 _2822_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net112),
    .B(_0831_),
    .A(_0830_),
    .Y(_0832_));
 sky130_as_sc_hs__mux2_2 _2823_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0597_),
    .B(_0832_),
    .A(_0829_),
    .Y(_0833_));
 sky130_as_sc_hs__ao22_2 _2824_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0607_),
    .C(_0833_),
    .B(_0826_),
    .D(_0610_),
    .Y(_0834_));
 sky130_as_sc_hs__or2_2 _2825_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net6),
    .B(_0643_),
    .Y(_0835_));
 sky130_as_sc_hs__oai21_2 _2826_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net24),
    .B(_0834_),
    .C(_0835_),
    .Y(_0836_));
 sky130_as_sc_hs__oa21_2 _2827_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net14),
    .B(_0640_),
    .C(_0587_),
    .Y(_0837_));
 sky130_as_sc_hs__aoi21_2 _2828_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\imm_buff[4] ),
    .B(net22),
    .C(_0837_),
    .Y(_0838_));
 sky130_as_sc_hs__ao31_2 _2829_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0787_),
    .B(_0819_),
    .C(_0836_),
    .D(_0838_),
    .Y(_0839_));
 sky130_as_sc_hs__clkbuff_4 _2830_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0839_),
    .Y(_0840_));
 sky130_as_sc_hs__inv_2 _2831_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_0840_),
    .Y(_0841_));
 sky130_as_sc_hs__buff_4 _2832_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0841_),
    .Y(_0842_));
 sky130_as_sc_hs__mux2_2 _2833_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0653_),
    .B(net50),
    .A(_0842_),
    .Y(_0843_));
 sky130_as_sc_hs__mux2_2 _2834_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0757_),
    .B(\last_MAR[4] ),
    .A(net50),
    .Y(_0844_));
 sky130_as_sc_hs__ao22_2 _2835_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0675_),
    .C(_0844_),
    .B(_0843_),
    .D(_0759_),
    .Y(_0845_));
 sky130_as_sc_hs__ao22_2 _2836_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net50),
    .C(_0845_),
    .B(_0665_),
    .D(_0761_),
    .Y(_0846_));
 sky130_as_sc_hs__mux2_2 _2837_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0672_),
    .B(_0846_),
    .A(\ROM_spi_dat_out[4] ),
    .Y(_0847_));
 sky130_as_sc_hs__and2_2 _2838_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net149),
    .B(_0847_),
    .Y(_0848_));
 sky130_as_sc_hs__buff_2 _2839_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0848_),
    .Y(_0004_));
 sky130_as_sc_hs__mux2_2 _2840_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net75),
    .B(\RAM[54][5] ),
    .A(\RAM[52][5] ),
    .Y(_0849_));
 sky130_as_sc_hs__mux2_2 _2841_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net75),
    .B(\RAM[55][5] ),
    .A(\RAM[53][5] ),
    .Y(_0850_));
 sky130_as_sc_hs__mux2_2 _2842_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net112),
    .B(_0850_),
    .A(_0849_),
    .Y(_0851_));
 sky130_as_sc_hs__mux2_2 _2843_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net67),
    .B(\RAM[50][5] ),
    .A(\RAM[48][5] ),
    .Y(_0852_));
 sky130_as_sc_hs__mux2_2 _2844_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net75),
    .B(\RAM[51][5] ),
    .A(\RAM[49][5] ),
    .Y(_0853_));
 sky130_as_sc_hs__mux2_2 _2845_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net112),
    .B(_0853_),
    .A(_0852_),
    .Y(_0854_));
 sky130_as_sc_hs__buff_6 _2846_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0597_),
    .Y(_0855_));
 sky130_as_sc_hs__mux2_2 _2847_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0855_),
    .B(_0854_),
    .A(_0851_),
    .Y(_0856_));
 sky130_as_sc_hs__mux2_2 _2848_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net81),
    .B(\RAM[62][5] ),
    .A(uo_out[5]),
    .Y(_0857_));
 sky130_as_sc_hs__mux2_2 _2849_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net81),
    .B(uio_out[5]),
    .A(\RAM[61][5] ),
    .Y(_0858_));
 sky130_as_sc_hs__mux2_2 _2850_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net117),
    .B(_0858_),
    .A(_0857_),
    .Y(_0859_));
 sky130_as_sc_hs__mux2_2 _2851_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net101),
    .B(\RAM[58][5] ),
    .A(\RAM[56][5] ),
    .Y(_0860_));
 sky130_as_sc_hs__mux2_2 _2852_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net78),
    .B(uio_oe[5]),
    .A(\RAM[57][5] ),
    .Y(_0861_));
 sky130_as_sc_hs__mux2_2 _2853_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net113),
    .B(_0861_),
    .A(_0860_),
    .Y(_0862_));
 sky130_as_sc_hs__mux2_2 _2854_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0855_),
    .B(_0862_),
    .A(_0859_),
    .Y(_0863_));
 sky130_as_sc_hs__mux2_2 _2855_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net55),
    .B(_0863_),
    .A(_0856_),
    .Y(_0864_));
 sky130_as_sc_hs__nor2_2 _2856_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0535_),
    .B(_0746_),
    .Y(_0865_));
 sky130_as_sc_hs__mux2_2 _2857_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net67),
    .B(\RAM[38][5] ),
    .A(\RAM[36][5] ),
    .Y(_0866_));
 sky130_as_sc_hs__mux2_2 _2858_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net67),
    .B(\RAM[39][5] ),
    .A(\RAM[37][5] ),
    .Y(_0867_));
 sky130_as_sc_hs__mux2_2 _2859_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net106),
    .B(_0867_),
    .A(_0866_),
    .Y(_0868_));
 sky130_as_sc_hs__mux2_2 _2860_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net64),
    .B(\RAM[34][5] ),
    .A(\RAM[32][5] ),
    .Y(_0869_));
 sky130_as_sc_hs__mux2_2 _2861_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net64),
    .B(\RAM[35][5] ),
    .A(\RAM[33][5] ),
    .Y(_0870_));
 sky130_as_sc_hs__mux2_2 _2862_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net104),
    .B(_0870_),
    .A(_0869_),
    .Y(_0871_));
 sky130_as_sc_hs__mux2_2 _2863_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0855_),
    .B(_0871_),
    .A(_0868_),
    .Y(_0872_));
 sky130_as_sc_hs__mux2_2 _2864_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net78),
    .B(\RAM[46][5] ),
    .A(\RAM[44][5] ),
    .Y(_0873_));
 sky130_as_sc_hs__mux2_2 _2865_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net79),
    .B(\RAM[47][5] ),
    .A(\RAM[45][5] ),
    .Y(_0874_));
 sky130_as_sc_hs__mux2_2 _2866_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net113),
    .B(_0874_),
    .A(_0873_),
    .Y(_0875_));
 sky130_as_sc_hs__mux2_2 _2867_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net76),
    .B(\RAM[42][5] ),
    .A(\RAM[40][5] ),
    .Y(_0876_));
 sky130_as_sc_hs__mux2_2 _2868_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net76),
    .B(\RAM[43][5] ),
    .A(\RAM[41][5] ),
    .Y(_0877_));
 sky130_as_sc_hs__mux2_2 _2869_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net112),
    .B(_0877_),
    .A(_0876_),
    .Y(_0878_));
 sky130_as_sc_hs__mux2_2 _2870_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0855_),
    .B(_0878_),
    .A(_0875_),
    .Y(_0879_));
 sky130_as_sc_hs__mux2_2 _2871_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net55),
    .B(_0879_),
    .A(_0872_),
    .Y(_0880_));
 sky130_as_sc_hs__ao22_2 _2872_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0864_),
    .C(_0880_),
    .B(_0865_),
    .D(_0535_),
    .Y(_0881_));
 sky130_as_sc_hs__ao21_2 _2873_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net7),
    .B(net24),
    .C(_0747_),
    .Y(_0882_));
 sky130_as_sc_hs__aoi21_2 _2874_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net140),
    .B(_0881_),
    .C(_0882_),
    .Y(_0883_));
 sky130_as_sc_hs__oai21_2 _2875_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net15),
    .B(_0640_),
    .C(_0587_),
    .Y(_0884_));
 sky130_as_sc_hs__inv_2 _2876_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\imm_buff[5] ),
    .Y(_0885_));
 sky130_as_sc_hs__mux2_2 _2877_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net72),
    .B(\RAM[22][5] ),
    .A(\RAM[20][5] ),
    .Y(_0886_));
 sky130_as_sc_hs__mux2_2 _2878_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net72),
    .B(\RAM[23][5] ),
    .A(\RAM[21][5] ),
    .Y(_0887_));
 sky130_as_sc_hs__mux2_2 _2879_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net110),
    .B(_0887_),
    .A(_0886_),
    .Y(_0888_));
 sky130_as_sc_hs__mux2_2 _2880_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net65),
    .B(\RAM[18][5] ),
    .A(\RAM[16][5] ),
    .Y(_0889_));
 sky130_as_sc_hs__mux2_2 _2881_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net65),
    .B(\RAM[19][5] ),
    .A(\RAM[17][5] ),
    .Y(_0890_));
 sky130_as_sc_hs__mux2_2 _2882_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net104),
    .B(_0890_),
    .A(_0889_),
    .Y(_0891_));
 sky130_as_sc_hs__mux2_2 _2883_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0855_),
    .B(_0891_),
    .A(_0888_),
    .Y(_0892_));
 sky130_as_sc_hs__mux2_2 _2884_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net71),
    .B(\RAM[30][5] ),
    .A(\RAM[28][5] ),
    .Y(_0893_));
 sky130_as_sc_hs__mux2_2 _2885_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net71),
    .B(\RAM[31][5] ),
    .A(\RAM[29][5] ),
    .Y(_0894_));
 sky130_as_sc_hs__mux2_2 _2886_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net109),
    .B(_0894_),
    .A(_0893_),
    .Y(_0895_));
 sky130_as_sc_hs__mux2_2 _2887_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net97),
    .B(\RAM[26][5] ),
    .A(\RAM[24][5] ),
    .Y(_0896_));
 sky130_as_sc_hs__mux2_2 _2888_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net97),
    .B(\RAM[27][5] ),
    .A(\RAM[25][5] ),
    .Y(_0897_));
 sky130_as_sc_hs__mux2_2 _2889_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net120),
    .B(_0897_),
    .A(_0896_),
    .Y(_0898_));
 sky130_as_sc_hs__mux2_2 _2890_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0855_),
    .B(_0898_),
    .A(_0895_),
    .Y(_0899_));
 sky130_as_sc_hs__ao22_2 _2891_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0562_),
    .C(_0899_),
    .B(_0892_),
    .D(_0553_),
    .Y(_0900_));
 sky130_as_sc_hs__mux2_2 _2892_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net66),
    .B(\RAM[3][5] ),
    .A(\RAM[1][5] ),
    .Y(_0901_));
 sky130_as_sc_hs__mux2_2 _2893_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net71),
    .B(\RAM[7][5] ),
    .A(\RAM[5][5] ),
    .Y(_0902_));
 sky130_as_sc_hs__mux2_2 _2894_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net56),
    .B(_0902_),
    .A(_0901_),
    .Y(_0903_));
 sky130_as_sc_hs__mux2_2 _2895_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net70),
    .B(\RAM[2][5] ),
    .A(\RAM[0][5] ),
    .Y(_0904_));
 sky130_as_sc_hs__mux2_2 _2896_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net70),
    .B(\RAM[6][5] ),
    .A(\RAM[4][5] ),
    .Y(_0905_));
 sky130_as_sc_hs__mux2_2 _2897_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net56),
    .B(_0905_),
    .A(_0904_),
    .Y(_0906_));
 sky130_as_sc_hs__mux2_2 _2898_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0620_),
    .B(_0906_),
    .A(_0903_),
    .Y(_0907_));
 sky130_as_sc_hs__mux2_2 _2899_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net99),
    .B(\RAM[14][5] ),
    .A(\RAM[12][5] ),
    .Y(_0908_));
 sky130_as_sc_hs__mux2_2 _2900_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net99),
    .B(\RAM[15][5] ),
    .A(\RAM[13][5] ),
    .Y(_0909_));
 sky130_as_sc_hs__mux2_2 _2901_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net120),
    .B(_0909_),
    .A(_0908_),
    .Y(_0910_));
 sky130_as_sc_hs__mux2_2 _2902_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net98),
    .B(\RAM[10][5] ),
    .A(\RAM[8][5] ),
    .Y(_0911_));
 sky130_as_sc_hs__mux2_2 _2903_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net98),
    .B(\RAM[11][5] ),
    .A(\RAM[9][5] ),
    .Y(_0912_));
 sky130_as_sc_hs__mux2_2 _2904_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net120),
    .B(_0912_),
    .A(_0911_),
    .Y(_0913_));
 sky130_as_sc_hs__mux2_2 _2905_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0855_),
    .B(_0913_),
    .A(_0910_),
    .Y(_0914_));
 sky130_as_sc_hs__oa22_2 _2906_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0589_),
    .B(_0907_),
    .C(_0914_),
    .D(_0631_),
    .Y(_0915_));
 sky130_as_sc_hs__iao211_2 _2907_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0788_),
    .B(_0900_),
    .C(_0915_),
    .D(_0635_),
    .Y(_0916_));
 sky130_as_sc_hs__mux2_2 _2908_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0587_),
    .B(_0916_),
    .A(_0885_),
    .Y(_0917_));
 sky130_as_sc_hs__oai21_2 _2909_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0883_),
    .B(_0884_),
    .C(_0917_),
    .Y(_0918_));
 sky130_as_sc_hs__mux2_2 _2910_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0653_),
    .B(net140),
    .A(_0918_),
    .Y(_0919_));
 sky130_as_sc_hs__buff_4 _2911_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0659_),
    .Y(_0920_));
 sky130_as_sc_hs__mux2_2 _2912_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0920_),
    .B(\last_MAR[5] ),
    .A(net140),
    .Y(_0921_));
 sky130_as_sc_hs__ao22_2 _2913_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0675_),
    .C(_0921_),
    .B(_0919_),
    .D(_0759_),
    .Y(_0922_));
 sky130_as_sc_hs__ao22_2 _2914_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net142),
    .C(_0922_),
    .B(_0665_),
    .D(_0761_),
    .Y(_0923_));
 sky130_as_sc_hs__mux2_2 _2915_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0672_),
    .B(_0923_),
    .A(\ROM_spi_dat_out[5] ),
    .Y(_0924_));
 sky130_as_sc_hs__and2_2 _2916_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net149),
    .B(_0924_),
    .Y(_0925_));
 sky130_as_sc_hs__buff_2 _2917_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0925_),
    .Y(_0005_));
 sky130_as_sc_hs__buff_2 _2918_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0534_),
    .Y(_0926_));
 sky130_as_sc_hs__or2_2 _2919_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net10),
    .B(_0640_),
    .Y(_0927_));
 sky130_as_sc_hs__and2_2 _2920_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net23),
    .B(_0927_),
    .Y(_0928_));
 sky130_as_sc_hs__mux2_2 _2921_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net77),
    .B(\RAM[42][0] ),
    .A(\RAM[40][0] ),
    .Y(_0929_));
 sky130_as_sc_hs__mux2_2 _2922_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net78),
    .B(\RAM[46][0] ),
    .A(\RAM[44][0] ),
    .Y(_0930_));
 sky130_as_sc_hs__mux2_2 _2923_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net60),
    .B(_0930_),
    .A(_0929_),
    .Y(_0931_));
 sky130_as_sc_hs__mux2_2 _2924_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net84),
    .B(\RAM[43][0] ),
    .A(\RAM[41][0] ),
    .Y(_0932_));
 sky130_as_sc_hs__ao21_2 _2925_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0698_),
    .B(_0932_),
    .C(_0630_),
    .Y(_0933_));
 sky130_as_sc_hs__mux2_2 _2926_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net88),
    .B(\RAM[47][0] ),
    .A(\RAM[45][0] ),
    .Y(_0934_));
 sky130_as_sc_hs__and2_2 _2927_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0695_),
    .B(_0934_),
    .Y(_0935_));
 sky130_as_sc_hs__aoi211_2 _2928_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_0931_),
    .C(_0933_),
    .D(_0935_),
    .Y(_0936_),
    .A(_0620_));
 sky130_as_sc_hs__mux2_2 _2929_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net87),
    .B(uio_oe[0]),
    .A(\RAM[57][0] ),
    .Y(_0937_));
 sky130_as_sc_hs__mux2_2 _2930_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net87),
    .B(\RAM[62][0] ),
    .A(uo_out[0]),
    .Y(_0938_));
 sky130_as_sc_hs__aoi22_2 _2931_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0698_),
    .B(_0937_),
    .C(_0938_),
    .D(_0700_),
    .Y(_0939_));
 sky130_as_sc_hs__mux2_2 _2932_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net101),
    .B(\RAM[58][0] ),
    .A(\RAM[56][0] ),
    .Y(_0940_));
 sky130_as_sc_hs__mux2_2 _2933_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net87),
    .B(uio_out[0]),
    .A(\RAM[61][0] ),
    .Y(_0941_));
 sky130_as_sc_hs__aoi22_2 _2934_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0703_),
    .B(_0940_),
    .C(_0941_),
    .D(_0694_),
    .Y(_0942_));
 sky130_as_sc_hs__ao31_2 _2935_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0641_),
    .B(_0939_),
    .C(_0942_),
    .D(_0737_),
    .Y(_0943_));
 sky130_as_sc_hs__or2_2 _2936_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0936_),
    .B(_0943_),
    .Y(_0944_));
 sky130_as_sc_hs__mux2_2 _2937_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net72),
    .B(\RAM[50][0] ),
    .A(\RAM[48][0] ),
    .Y(_0945_));
 sky130_as_sc_hs__mux2_2 _2938_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net85),
    .B(\RAM[51][0] ),
    .A(\RAM[49][0] ),
    .Y(_0946_));
 sky130_as_sc_hs__mux2_2 _2939_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net114),
    .B(_0946_),
    .A(_0945_),
    .Y(_0947_));
 sky130_as_sc_hs__mux2_2 _2940_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net85),
    .B(\RAM[54][0] ),
    .A(\RAM[52][0] ),
    .Y(_0948_));
 sky130_as_sc_hs__mux2_2 _2941_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net77),
    .B(\RAM[55][0] ),
    .A(\RAM[53][0] ),
    .Y(_0949_));
 sky130_as_sc_hs__mux2_2 _2942_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net115),
    .B(_0949_),
    .A(_0948_),
    .Y(_0950_));
 sky130_as_sc_hs__ao31_2 _2943_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net49),
    .B(net58),
    .C(_0950_),
    .D(net52),
    .Y(_0951_));
 sky130_as_sc_hs__mux2_2 _2944_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net72),
    .B(\RAM[38][0] ),
    .A(\RAM[36][0] ),
    .Y(_0952_));
 sky130_as_sc_hs__mux2_2 _2945_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net73),
    .B(\RAM[39][0] ),
    .A(\RAM[37][0] ),
    .Y(_0953_));
 sky130_as_sc_hs__mux2_2 _2946_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net110),
    .B(_0953_),
    .A(_0952_),
    .Y(_0954_));
 sky130_as_sc_hs__mux2_2 _2947_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net69),
    .B(\RAM[34][0] ),
    .A(\RAM[32][0] ),
    .Y(_0955_));
 sky130_as_sc_hs__mux2_2 _2948_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net64),
    .B(\RAM[35][0] ),
    .A(\RAM[33][0] ),
    .Y(_0956_));
 sky130_as_sc_hs__mux2_2 _2949_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net104),
    .B(_0956_),
    .A(_0955_),
    .Y(_0957_));
 sky130_as_sc_hs__ao22_2 _2950_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0684_),
    .C(_0957_),
    .B(_0954_),
    .D(_0683_),
    .Y(_0958_));
 sky130_as_sc_hs__aoi211_2 _2951_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_0947_),
    .C(_0951_),
    .D(_0958_),
    .Y(_0959_),
    .A(_0679_));
 sky130_as_sc_hs__aoi21_2 _2952_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net2),
    .B(net24),
    .C(_0747_),
    .Y(_0960_));
 sky130_as_sc_hs__mux2_2 _2953_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net90),
    .B(\RAM[31][0] ),
    .A(\RAM[29][0] ),
    .Y(_0961_));
 sky130_as_sc_hs__mux2_2 _2954_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net96),
    .B(\RAM[26][0] ),
    .A(\RAM[24][0] ),
    .Y(_0962_));
 sky130_as_sc_hs__aoi22_2 _2955_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0695_),
    .B(_0961_),
    .C(_0962_),
    .D(_0703_),
    .Y(_0963_));
 sky130_as_sc_hs__mux2_2 _2956_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net96),
    .B(\RAM[27][0] ),
    .A(\RAM[25][0] ),
    .Y(_0964_));
 sky130_as_sc_hs__mux2_2 _2957_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net90),
    .B(\RAM[30][0] ),
    .A(\RAM[28][0] ),
    .Y(_0965_));
 sky130_as_sc_hs__aoi22_2 _2958_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net26),
    .B(_0964_),
    .C(_0965_),
    .D(net25),
    .Y(_0966_));
 sky130_as_sc_hs__nand3_2 _2959_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0641_),
    .B(_0963_),
    .C(_0966_),
    .Y(_0967_));
 sky130_as_sc_hs__nor2_2 _2960_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0552_),
    .B(net51),
    .Y(_0968_));
 sky130_as_sc_hs__mux2_2 _2961_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net94),
    .B(\RAM[11][0] ),
    .A(\RAM[9][0] ),
    .Y(_0969_));
 sky130_as_sc_hs__mux2_2 _2962_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net96),
    .B(\RAM[10][0] ),
    .A(\RAM[8][0] ),
    .Y(_0970_));
 sky130_as_sc_hs__aoi22_2 _2963_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net26),
    .B(_0969_),
    .C(_0970_),
    .D(_0703_),
    .Y(_0971_));
 sky130_as_sc_hs__mux2_2 _2964_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net94),
    .B(\RAM[14][0] ),
    .A(\RAM[12][0] ),
    .Y(_0972_));
 sky130_as_sc_hs__mux2_2 _2965_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net93),
    .B(\RAM[15][0] ),
    .A(\RAM[13][0] ),
    .Y(_0973_));
 sky130_as_sc_hs__aoi22_2 _2966_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net25),
    .B(_0972_),
    .C(_0973_),
    .D(_0695_),
    .Y(_0974_));
 sky130_as_sc_hs__aoi31_2 _2967_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0968_),
    .B(_0971_),
    .C(_0974_),
    .D(net141),
    .Y(_0975_));
 sky130_as_sc_hs__nor2_2 _2968_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net54),
    .B(net51),
    .Y(_0976_));
 sky130_as_sc_hs__nand2_2 _2969_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0560_),
    .B(_0976_),
    .Y(_0977_));
 sky130_as_sc_hs__mux2_2 _2970_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net70),
    .B(\RAM[2][0] ),
    .A(\RAM[0][0] ),
    .Y(_0978_));
 sky130_as_sc_hs__mux2_2 _2971_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net71),
    .B(\RAM[3][0] ),
    .A(\RAM[1][0] ),
    .Y(_0979_));
 sky130_as_sc_hs__mux2_2 _2972_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net109),
    .B(_0979_),
    .A(_0978_),
    .Y(_0980_));
 sky130_as_sc_hs__nand2_2 _2973_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net62),
    .B(_0976_),
    .Y(_0981_));
 sky130_as_sc_hs__mux2_2 _2974_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net92),
    .B(\RAM[6][0] ),
    .A(\RAM[4][0] ),
    .Y(_0982_));
 sky130_as_sc_hs__mux2_2 _2975_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net92),
    .B(\RAM[7][0] ),
    .A(\RAM[5][0] ),
    .Y(_0983_));
 sky130_as_sc_hs__mux2_2 _2976_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net119),
    .B(_0983_),
    .A(_0982_),
    .Y(_0984_));
 sky130_as_sc_hs__oa22_2 _2977_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0977_),
    .B(_0980_),
    .C(_0981_),
    .D(_0984_),
    .Y(_0985_));
 sky130_as_sc_hs__mux2_2 _2978_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net67),
    .B(\RAM[18][0] ),
    .A(\RAM[16][0] ),
    .Y(_0986_));
 sky130_as_sc_hs__mux2_2 _2979_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net67),
    .B(\RAM[19][0] ),
    .A(\RAM[17][0] ),
    .Y(_0987_));
 sky130_as_sc_hs__mux2_2 _2980_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net106),
    .B(_0987_),
    .A(_0986_),
    .Y(_0988_));
 sky130_as_sc_hs__nor2b_2 _2981_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net52),
    .Y(_0989_),
    .B(net49));
 sky130_as_sc_hs__nand2_2 _2982_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0560_),
    .B(_0989_),
    .Y(_0990_));
 sky130_as_sc_hs__nand2_2 _2983_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net61),
    .B(_0989_),
    .Y(_0991_));
 sky130_as_sc_hs__mux2_2 _2984_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net93),
    .B(\RAM[22][0] ),
    .A(\RAM[20][0] ),
    .Y(_0992_));
 sky130_as_sc_hs__mux2_2 _2985_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net93),
    .B(\RAM[23][0] ),
    .A(\RAM[21][0] ),
    .Y(_0993_));
 sky130_as_sc_hs__mux2_2 _2986_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net119),
    .B(_0993_),
    .A(_0992_),
    .Y(_0994_));
 sky130_as_sc_hs__oa22_2 _2987_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0988_),
    .B(_0990_),
    .C(_0991_),
    .D(_0994_),
    .Y(_0995_));
 sky130_as_sc_hs__nand4_2 _2988_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0967_),
    .B(_0975_),
    .C(_0985_),
    .Y(_0996_),
    .D(_0995_));
 sky130_as_sc_hs__iao211_2 _2989_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0944_),
    .B(_0959_),
    .C(_0960_),
    .D(_0996_),
    .Y(_0997_));
 sky130_as_sc_hs__and2_2 _2990_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\imm_buff[0] ),
    .B(_0785_),
    .Y(_0998_));
 sky130_as_sc_hs__ao21_4 _2991_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0928_),
    .B(_0997_),
    .C(_0998_),
    .Y(_0999_));
 sky130_as_sc_hs__nor2_2 _2992_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net39),
    .B(net35),
    .Y(_1000_));
 sky130_as_sc_hs__nor2_2 _2993_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net45),
    .B(net41),
    .Y(_1001_));
 sky130_as_sc_hs__nand2_2 _2994_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1000_),
    .B(_1001_),
    .Y(_1002_));
 sky130_as_sc_hs__nand2_2 _2995_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\instr_cycle[1] ),
    .B(net33),
    .Y(_1003_));
 sky130_as_sc_hs__nor2_4 _2996_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1002_),
    .B(_1003_),
    .Y(_1004_));
 sky130_as_sc_hs__mux2_2 _2997_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1004_),
    .B(_0999_),
    .A(\P[0] ),
    .Y(_1005_));
 sky130_as_sc_hs__mux2_2 _2998_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0920_),
    .B(\last_P[0] ),
    .A(\P[0] ),
    .Y(_1006_));
 sky130_as_sc_hs__ao22_2 _2999_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0926_),
    .C(_1006_),
    .B(_1005_),
    .D(_0759_),
    .Y(_1007_));
 sky130_as_sc_hs__buff_2 _3000_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0533_),
    .Y(_1008_));
 sky130_as_sc_hs__ao22_2 _3001_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[0] ),
    .C(_1007_),
    .B(_0665_),
    .D(_1008_),
    .Y(_1009_));
 sky130_as_sc_hs__inv_2 _3002_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\ROM_dest[1] ),
    .Y(_1010_));
 sky130_as_sc_hs__nor2_2 _3003_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\ROM_dest[2] ),
    .B(_0670_),
    .Y(_1011_));
 sky130_as_sc_hs__nand2_4 _3004_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1010_),
    .B(_1011_),
    .Y(_1012_));
 sky130_as_sc_hs__mux2_2 _3005_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1012_),
    .B(_1009_),
    .A(\ROM_spi_dat_out[0] ),
    .Y(_1013_));
 sky130_as_sc_hs__and2_2 _3006_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net152),
    .B(_1013_),
    .Y(_1014_));
 sky130_as_sc_hs__buff_2 _3007_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1014_),
    .Y(_0006_));
 sky130_as_sc_hs__oai22_2 _3008_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net11),
    .B(_0640_),
    .C(_0643_),
    .D(net3),
    .Y(_1015_));
 sky130_as_sc_hs__nor2_4 _3009_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net22),
    .B(_1015_),
    .Y(_1016_));
 sky130_as_sc_hs__mux2_2 _3010_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net90),
    .B(\RAM[30][1] ),
    .A(\RAM[28][1] ),
    .Y(_1017_));
 sky130_as_sc_hs__mux2_2 _3011_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net92),
    .B(\RAM[31][1] ),
    .A(\RAM[29][1] ),
    .Y(_1018_));
 sky130_as_sc_hs__mux2_2 _3012_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net119),
    .B(_1018_),
    .A(_1017_),
    .Y(_1019_));
 sky130_as_sc_hs__mux2_2 _3013_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net97),
    .B(\RAM[26][1] ),
    .A(\RAM[24][1] ),
    .Y(_1020_));
 sky130_as_sc_hs__mux2_2 _3014_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net97),
    .B(\RAM[27][1] ),
    .A(\RAM[25][1] ),
    .Y(_1021_));
 sky130_as_sc_hs__mux2_2 _3015_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net120),
    .B(_1021_),
    .A(_1020_),
    .Y(_1022_));
 sky130_as_sc_hs__mux2_2 _3016_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0542_),
    .B(_1022_),
    .A(_1019_),
    .Y(_1023_));
 sky130_as_sc_hs__mux2_2 _3017_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net111),
    .B(\RAM[23][1] ),
    .A(\RAM[22][1] ),
    .Y(_1024_));
 sky130_as_sc_hs__or2_2 _3018_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0568_),
    .B(_1024_),
    .Y(_1025_));
 sky130_as_sc_hs__mux2_2 _3019_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net107),
    .B(\RAM[17][1] ),
    .A(\RAM[16][1] ),
    .Y(_1026_));
 sky130_as_sc_hs__mux2_2 _3020_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net106),
    .B(\RAM[19][1] ),
    .A(\RAM[18][1] ),
    .Y(_1027_));
 sky130_as_sc_hs__oa22_2 _3021_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0563_),
    .B(_1026_),
    .C(_1027_),
    .D(_0565_),
    .Y(_1028_));
 sky130_as_sc_hs__mux2_2 _3022_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net110),
    .B(\RAM[21][1] ),
    .A(\RAM[20][1] ),
    .Y(_1029_));
 sky130_as_sc_hs__oa21_2 _3023_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0571_),
    .B(_1029_),
    .C(_0562_),
    .Y(_1030_));
 sky130_as_sc_hs__ao31_2 _3024_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1025_),
    .B(_1028_),
    .C(_1030_),
    .D(_0788_),
    .Y(_1031_));
 sky130_as_sc_hs__ao21_2 _3025_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0553_),
    .B(_1023_),
    .C(_1031_),
    .Y(_1032_));
 sky130_as_sc_hs__mux2_2 _3026_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net97),
    .B(\RAM[10][1] ),
    .A(\RAM[8][1] ),
    .Y(_1033_));
 sky130_as_sc_hs__mux2_2 _3027_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net98),
    .B(\RAM[14][1] ),
    .A(\RAM[12][1] ),
    .Y(_1034_));
 sky130_as_sc_hs__mux2_2 _3028_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net62),
    .B(_1034_),
    .A(_1033_),
    .Y(_1035_));
 sky130_as_sc_hs__nor3_2 _3029_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net121),
    .B(_0631_),
    .C(_1035_),
    .Y(_1036_));
 sky130_as_sc_hs__mux2_2 _3030_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net99),
    .B(\RAM[11][1] ),
    .A(\RAM[9][1] ),
    .Y(_1037_));
 sky130_as_sc_hs__mux2_2 _3031_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net99),
    .B(\RAM[15][1] ),
    .A(\RAM[13][1] ),
    .Y(_1038_));
 sky130_as_sc_hs__mux2_2 _3032_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net62),
    .B(_1038_),
    .A(_1037_),
    .Y(_1039_));
 sky130_as_sc_hs__nor3_2 _3033_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0620_),
    .B(_0631_),
    .C(_1039_),
    .Y(_1040_));
 sky130_as_sc_hs__mux2_2 _3034_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net92),
    .B(\RAM[6][1] ),
    .A(\RAM[4][1] ),
    .Y(_1041_));
 sky130_as_sc_hs__mux2_2 _3035_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net92),
    .B(\RAM[7][1] ),
    .A(\RAM[5][1] ),
    .Y(_1042_));
 sky130_as_sc_hs__mux2_2 _3036_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net119),
    .B(_1042_),
    .A(_1041_),
    .Y(_1043_));
 sky130_as_sc_hs__mux2_2 _3037_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net70),
    .B(\RAM[2][1] ),
    .A(\RAM[0][1] ),
    .Y(_1044_));
 sky130_as_sc_hs__mux2_2 _3038_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net70),
    .B(\RAM[3][1] ),
    .A(\RAM[1][1] ),
    .Y(_1045_));
 sky130_as_sc_hs__mux2_2 _3039_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net109),
    .B(_1045_),
    .A(_1044_),
    .Y(_1046_));
 sky130_as_sc_hs__oai22_2 _3040_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0981_),
    .B(_1043_),
    .C(_1046_),
    .D(_0977_),
    .Y(_1047_));
 sky130_as_sc_hs__nor3_2 _3041_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1036_),
    .B(_1040_),
    .C(_1047_),
    .Y(_1048_));
 sky130_as_sc_hs__mux2_2 _3042_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net84),
    .B(\RAM[58][1] ),
    .A(\RAM[56][1] ),
    .Y(_1049_));
 sky130_as_sc_hs__or2_2 _3043_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0625_),
    .B(_1049_),
    .Y(_1050_));
 sky130_as_sc_hs__inv_2 _3044_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\RAM[62][1] ),
    .Y(_1051_));
 sky130_as_sc_hs__aoi31_2 _3045_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net84),
    .B(_1051_),
    .C(_0700_),
    .D(_0638_),
    .Y(_1052_));
 sky130_as_sc_hs__nand2_2 _3046_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net115),
    .B(net59),
    .Y(_1053_));
 sky130_as_sc_hs__mux2_2 _3047_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net87),
    .B(uio_out[1]),
    .A(\RAM[61][1] ),
    .Y(_1054_));
 sky130_as_sc_hs__mux2_2 _3048_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net86),
    .B(uio_oe[1]),
    .A(\RAM[57][1] ),
    .Y(_1055_));
 sky130_as_sc_hs__nand2b_2 _3049_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(net114),
    .Y(_1056_),
    .A(net59));
 sky130_as_sc_hs__oa22_2 _3050_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1053_),
    .B(_1054_),
    .C(_1055_),
    .D(_1056_),
    .Y(_1057_));
 sky130_as_sc_hs__nand3_2 _3051_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1050_),
    .B(_1052_),
    .C(_1057_),
    .Y(_1058_));
 sky130_as_sc_hs__mux2_2 _3052_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net85),
    .B(\RAM[42][1] ),
    .A(\RAM[40][1] ),
    .Y(_1059_));
 sky130_as_sc_hs__mux2_2 _3053_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net86),
    .B(\RAM[46][1] ),
    .A(\RAM[44][1] ),
    .Y(_1060_));
 sky130_as_sc_hs__oa22_2 _3054_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0625_),
    .B(_1059_),
    .C(_1060_),
    .D(_0627_),
    .Y(_1061_));
 sky130_as_sc_hs__mux2_2 _3055_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net86),
    .B(\RAM[43][1] ),
    .A(\RAM[41][1] ),
    .Y(_1062_));
 sky130_as_sc_hs__mux2_2 _3056_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net87),
    .B(\RAM[47][1] ),
    .A(\RAM[45][1] ),
    .Y(_1063_));
 sky130_as_sc_hs__oa22_2 _3057_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1056_),
    .B(_1062_),
    .C(_1063_),
    .D(_1053_),
    .Y(_1064_));
 sky130_as_sc_hs__nand3_2 _3058_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0632_),
    .B(_1061_),
    .C(_1064_),
    .Y(_1065_));
 sky130_as_sc_hs__mux2_2 _3059_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net110),
    .B(\RAM[37][1] ),
    .A(\RAM[36][1] ),
    .Y(_1066_));
 sky130_as_sc_hs__mux2_2 _3060_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net110),
    .B(\RAM[39][1] ),
    .A(\RAM[38][1] ),
    .Y(_1067_));
 sky130_as_sc_hs__oa22_2 _3061_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0571_),
    .B(_1066_),
    .C(_1067_),
    .D(_0568_),
    .Y(_1068_));
 sky130_as_sc_hs__mux2_2 _3062_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net105),
    .B(\RAM[35][1] ),
    .A(\RAM[34][1] ),
    .Y(_1069_));
 sky130_as_sc_hs__mux2_2 _3063_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net104),
    .B(\RAM[33][1] ),
    .A(\RAM[32][1] ),
    .Y(_1070_));
 sky130_as_sc_hs__oa22_2 _3064_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0565_),
    .B(_1069_),
    .C(_1070_),
    .D(_0563_),
    .Y(_1071_));
 sky130_as_sc_hs__nand3_2 _3065_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0590_),
    .B(_1068_),
    .C(_1071_),
    .Y(_1072_));
 sky130_as_sc_hs__mux2_2 _3066_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net85),
    .B(\RAM[51][1] ),
    .A(\RAM[49][1] ),
    .Y(_1073_));
 sky130_as_sc_hs__mux2_2 _3067_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net84),
    .B(\RAM[50][1] ),
    .A(\RAM[48][1] ),
    .Y(_1074_));
 sky130_as_sc_hs__oa22_2 _3068_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1056_),
    .B(_1073_),
    .C(_1074_),
    .D(_0625_),
    .Y(_1075_));
 sky130_as_sc_hs__mux2_2 _3069_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net85),
    .B(\RAM[54][1] ),
    .A(\RAM[52][1] ),
    .Y(_1076_));
 sky130_as_sc_hs__mux2_2 _3070_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net85),
    .B(\RAM[55][1] ),
    .A(\RAM[53][1] ),
    .Y(_1077_));
 sky130_as_sc_hs__oa22_2 _3071_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0627_),
    .B(_1076_),
    .C(_1077_),
    .D(_1053_),
    .Y(_1078_));
 sky130_as_sc_hs__aoi31_2 _3072_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0610_),
    .B(_1075_),
    .C(_1078_),
    .D(_0747_),
    .Y(_1079_));
 sky130_as_sc_hs__nand4_2 _3073_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1058_),
    .B(_1065_),
    .C(_1072_),
    .Y(_1080_),
    .D(_1079_));
 sky130_as_sc_hs__ao21_2 _3074_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1032_),
    .B(_1048_),
    .C(_1080_),
    .Y(_1081_));
 sky130_as_sc_hs__and2_2 _3075_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\imm_buff[1] ),
    .B(net22),
    .Y(_1082_));
 sky130_as_sc_hs__ao21_2 _3076_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1016_),
    .B(_1081_),
    .C(_1082_),
    .Y(_1083_));
 sky130_as_sc_hs__buff_4 _3077_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1083_),
    .Y(_1084_));
 sky130_as_sc_hs__mux2_2 _3078_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1004_),
    .B(_1084_),
    .A(\P[1] ),
    .Y(_1085_));
 sky130_as_sc_hs__mux2_2 _3079_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0920_),
    .B(\last_P[1] ),
    .A(\P[1] ),
    .Y(_1086_));
 sky130_as_sc_hs__ao22_2 _3080_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0926_),
    .C(_1086_),
    .B(_1085_),
    .D(_0759_),
    .Y(_1087_));
 sky130_as_sc_hs__ao22_2 _3081_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[1] ),
    .C(_1087_),
    .B(_0665_),
    .D(_1008_),
    .Y(_1088_));
 sky130_as_sc_hs__mux2_2 _3082_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1012_),
    .B(_1088_),
    .A(\ROM_spi_dat_out[1] ),
    .Y(_1089_));
 sky130_as_sc_hs__and2_2 _3083_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net152),
    .B(_1089_),
    .Y(_1090_));
 sky130_as_sc_hs__buff_2 _3084_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1090_),
    .Y(_0007_));
 sky130_as_sc_hs__buff_2 _3085_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0664_),
    .Y(_1091_));
 sky130_as_sc_hs__inv_2 _3086_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\P[2] ),
    .Y(_1092_));
 sky130_as_sc_hs__oai21_2 _3087_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0576_),
    .B(_0637_),
    .C(_0645_),
    .Y(_1093_));
 sky130_as_sc_hs__clkbuff_4 _3088_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1093_),
    .Y(_1094_));
 sky130_as_sc_hs__mux2_2 _3089_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1004_),
    .B(_1094_),
    .A(_1092_),
    .Y(_1095_));
 sky130_as_sc_hs__inv_2 _3090_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_1095_),
    .Y(_1096_));
 sky130_as_sc_hs__mux2_2 _3091_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0920_),
    .B(\last_P[2] ),
    .A(\P[2] ),
    .Y(_1097_));
 sky130_as_sc_hs__ao22_2 _3092_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0926_),
    .C(_1097_),
    .B(_1096_),
    .D(_0759_),
    .Y(_1098_));
 sky130_as_sc_hs__ao22_2 _3093_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[2] ),
    .C(_1098_),
    .B(_1091_),
    .D(_1008_),
    .Y(_1099_));
 sky130_as_sc_hs__mux2_2 _3094_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1012_),
    .B(_1099_),
    .A(\ROM_spi_dat_out[2] ),
    .Y(_1100_));
 sky130_as_sc_hs__and2_2 _3095_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net154),
    .B(_1100_),
    .Y(_1101_));
 sky130_as_sc_hs__buff_2 _3096_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1101_),
    .Y(_0008_));
 sky130_as_sc_hs__nor2_2 _3097_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\P[3] ),
    .B(_1004_),
    .Y(_1102_));
 sky130_as_sc_hs__aoi21_2 _3098_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0754_),
    .B(_1004_),
    .C(_1102_),
    .Y(_1103_));
 sky130_as_sc_hs__mux2_2 _3099_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0920_),
    .B(\last_P[3] ),
    .A(\P[3] ),
    .Y(_1104_));
 sky130_as_sc_hs__ao22_2 _3100_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0926_),
    .C(_1104_),
    .B(_1103_),
    .D(_0759_),
    .Y(_1105_));
 sky130_as_sc_hs__ao22_2 _3101_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[3] ),
    .C(_1105_),
    .B(_1091_),
    .D(_1008_),
    .Y(_1106_));
 sky130_as_sc_hs__mux2_2 _3102_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1012_),
    .B(_1106_),
    .A(\ROM_spi_dat_out[3] ),
    .Y(_1107_));
 sky130_as_sc_hs__and2_2 _3103_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net154),
    .B(_1107_),
    .Y(_1108_));
 sky130_as_sc_hs__buff_2 _3104_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1108_),
    .Y(_0009_));
 sky130_as_sc_hs__mux2_2 _3105_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1004_),
    .B(_0842_),
    .A(\P[4] ),
    .Y(_1109_));
 sky130_as_sc_hs__mux2_2 _3106_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0920_),
    .B(\last_P[4] ),
    .A(\P[4] ),
    .Y(_1110_));
 sky130_as_sc_hs__ao22_2 _3107_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0926_),
    .C(_1110_),
    .B(_1109_),
    .D(_0657_),
    .Y(_1111_));
 sky130_as_sc_hs__ao22_2 _3108_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[4] ),
    .C(_1111_),
    .B(_1091_),
    .D(_1008_),
    .Y(_1112_));
 sky130_as_sc_hs__mux2_2 _3109_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1012_),
    .B(_1112_),
    .A(\ROM_spi_dat_out[4] ),
    .Y(_1113_));
 sky130_as_sc_hs__and2_2 _3110_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net155),
    .B(_1113_),
    .Y(_1114_));
 sky130_as_sc_hs__buff_2 _3111_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1114_),
    .Y(_0010_));
 sky130_as_sc_hs__mux2_2 _3112_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1004_),
    .B(_0918_),
    .A(\P[5] ),
    .Y(_1115_));
 sky130_as_sc_hs__mux2_2 _3113_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0920_),
    .B(\last_P[5] ),
    .A(\P[5] ),
    .Y(_1116_));
 sky130_as_sc_hs__ao22_2 _3114_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0926_),
    .C(_1116_),
    .B(_1115_),
    .D(_0657_),
    .Y(_1117_));
 sky130_as_sc_hs__ao22_2 _3115_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[5] ),
    .C(_1117_),
    .B(_1091_),
    .D(_1008_),
    .Y(_1118_));
 sky130_as_sc_hs__mux2_2 _3116_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1012_),
    .B(_1118_),
    .A(\ROM_spi_dat_out[5] ),
    .Y(_1119_));
 sky130_as_sc_hs__and2_2 _3117_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net155),
    .B(_1119_),
    .Y(_1120_));
 sky130_as_sc_hs__buff_2 _3118_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1120_),
    .Y(_0011_));
 sky130_as_sc_hs__or2_2 _3119_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0655_),
    .B(_0659_),
    .Y(_1121_));
 sky130_as_sc_hs__nand2_2 _3120_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net28),
    .B(_1001_),
    .Y(_1122_));
 sky130_as_sc_hs__inv_2 _3121_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net45),
    .Y(_1123_));
 sky130_as_sc_hs__mux2_2 _3122_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net41),
    .B(net28),
    .A(_1123_),
    .Y(_1124_));
 sky130_as_sc_hs__mux2_2 _3123_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net32),
    .B(_1124_),
    .A(_1122_),
    .Y(_1125_));
 sky130_as_sc_hs__nor2_2 _3124_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0658_),
    .B(_1125_),
    .Y(_1126_));
 sky130_as_sc_hs__or2_2 _3125_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1121_),
    .B(_1126_),
    .Y(_1127_));
 sky130_as_sc_hs__clkbuff_4 _3126_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0648_),
    .Y(_1128_));
 sky130_as_sc_hs__clkbuff_4 _3127_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1128_),
    .Y(_1129_));
 sky130_as_sc_hs__inv_2 _3128_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net149),
    .Y(_1130_));
 sky130_as_sc_hs__ao31_2 _3129_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1129_),
    .B(_0578_),
    .C(_0652_),
    .D(_1130_),
    .Y(_1131_));
 sky130_as_sc_hs__nor3_2 _3130_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1091_),
    .B(_1127_),
    .C(_1131_),
    .Y(_1132_));
 sky130_as_sc_hs__nor2_2 _3131_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1123_),
    .B(_1128_),
    .Y(_1133_));
 sky130_as_sc_hs__inv_2 _3132_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_1133_),
    .Y(_1134_));
 sky130_as_sc_hs__oa21_2 _3133_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net34),
    .B(net40),
    .C(_0583_),
    .Y(_1135_));
 sky130_as_sc_hs__oa22_2 _3134_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1134_),
    .B(_0581_),
    .C(_1135_),
    .D(net29),
    .Y(_1136_));
 sky130_as_sc_hs__nor2_2 _3135_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0584_),
    .B(_1136_),
    .Y(_1137_));
 sky130_as_sc_hs__inv_2 _3136_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net32),
    .Y(_1138_));
 sky130_as_sc_hs__buff_4 _3137_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1138_),
    .Y(_1139_));
 sky130_as_sc_hs__oa21_2 _3138_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1139_),
    .B(_0580_),
    .C(net29),
    .Y(_1140_));
 sky130_as_sc_hs__or2_2 _3139_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net45),
    .B(net41),
    .Y(_1141_));
 sky130_as_sc_hs__mux2_2 _3140_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net33),
    .B(_1124_),
    .A(_1141_),
    .Y(_1142_));
 sky130_as_sc_hs__nor2_2 _3141_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0655_),
    .B(_0660_),
    .Y(_1143_));
 sky130_as_sc_hs__oai21_2 _3142_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0658_),
    .B(_1142_),
    .C(_1143_),
    .Y(_1144_));
 sky130_as_sc_hs__or2_2 _3143_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0530_),
    .B(_0532_),
    .Y(_1145_));
 sky130_as_sc_hs__buff_4 _3144_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1145_),
    .Y(_1146_));
 sky130_as_sc_hs__ao21_2 _3145_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0663_),
    .B(_1144_),
    .C(_1146_),
    .Y(_1147_));
 sky130_as_sc_hs__ao22_2 _3146_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1132_),
    .C(_1147_),
    .B(_1140_),
    .D(net160),
    .Y(_1148_));
 sky130_as_sc_hs__ao22_2 _3147_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1132_),
    .C(_1148_),
    .B(_1137_),
    .D(\ROM_dest[1] ),
    .Y(_1149_));
 sky130_as_sc_hs__buff_2 _3148_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1149_),
    .Y(_0019_));
 sky130_as_sc_hs__inv_4 _3149_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net37),
    .Y(_1150_));
 sky130_as_sc_hs__clkbuff_4 _3150_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1150_),
    .Y(_1151_));
 sky130_as_sc_hs__nor2_2 _3151_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net45),
    .B(_0577_),
    .Y(_1152_));
 sky130_as_sc_hs__aoi31_2 _3152_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1151_),
    .B(net33),
    .C(_1152_),
    .D(net28),
    .Y(_1153_));
 sky130_as_sc_hs__oa21_2 _3153_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0584_),
    .B(_1135_),
    .C(_1153_),
    .Y(_1154_));
 sky130_as_sc_hs__ao22_2 _3154_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_dest[2] ),
    .C(_1154_),
    .B(_1148_),
    .D(_1132_),
    .Y(_1155_));
 sky130_as_sc_hs__buff_2 _3155_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1155_),
    .Y(_0020_));
 sky130_as_sc_hs__buff_4 _3156_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1130_),
    .Y(_1156_));
 sky130_as_sc_hs__buff_8 _3157_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1156_),
    .Y(_1157_));
 sky130_as_sc_hs__buff_8 _3158_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1157_),
    .Y(_1158_));
 sky130_as_sc_hs__buff_4 _3159_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0656_),
    .Y(_1159_));
 sky130_as_sc_hs__mux2_2 _3160_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1146_),
    .B(_1159_),
    .A(_0663_),
    .Y(_1160_));
 sky130_as_sc_hs__nor2_2 _3161_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1158_),
    .B(_1160_),
    .Y(_0023_));
 sky130_as_sc_hs__nor2_2 _3162_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1121_),
    .B(_1126_),
    .Y(_1161_));
 sky130_as_sc_hs__nor2_2 _3163_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0648_),
    .B(_0783_),
    .Y(_1162_));
 sky130_as_sc_hs__nand4_2 _3164_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net37),
    .B(_1139_),
    .C(net45),
    .Y(_1163_),
    .D(_1162_));
 sky130_as_sc_hs__ao21_2 _3165_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1002_),
    .B(_1163_),
    .C(net28),
    .Y(_1164_));
 sky130_as_sc_hs__nand3_2 _3166_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0761_),
    .B(_1161_),
    .C(_1164_),
    .Y(_1165_));
 sky130_as_sc_hs__nand2_2 _3167_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net594),
    .B(_1146_),
    .Y(_1166_));
 sky130_as_sc_hs__aoi21_2 _3168_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1165_),
    .B(_1166_),
    .C(_1158_),
    .Y(_0022_));
 sky130_as_sc_hs__nor2_2 _3169_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net139),
    .B(_0761_),
    .Y(_1167_));
 sky130_as_sc_hs__nand2_2 _3170_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net32),
    .B(_1000_),
    .Y(_1168_));
 sky130_as_sc_hs__inv_2 _3171_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net30),
    .Y(_1169_));
 sky130_as_sc_hs__aoi21_2 _3172_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1134_),
    .B(_1141_),
    .C(_1169_),
    .Y(_1170_));
 sky130_as_sc_hs__oa21_2 _3173_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net28),
    .B(_0580_),
    .C(_1002_),
    .Y(_1171_));
 sky130_as_sc_hs__oai22_2 _3174_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1168_),
    .B(_1170_),
    .C(_1171_),
    .D(net32),
    .Y(_1172_));
 sky130_as_sc_hs__aoi211_2 _3175_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1172_),
    .C(_1146_),
    .D(net590),
    .Y(_1173_),
    .A(net136));
 sky130_as_sc_hs__oai21_2 _3176_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1167_),
    .B(_1173_),
    .C(net160),
    .Y(_0021_));
 sky130_as_sc_hs__nand2_2 _3177_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net168),
    .B(_1148_),
    .Y(_1174_));
 sky130_as_sc_hs__iao211_2 _3178_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0663_),
    .B(_1146_),
    .C(_1174_),
    .D(net157),
    .Y(_0018_));
 sky130_as_sc_hs__inv_2 _3179_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\RAM[58][2] ),
    .Y(_1175_));
 sky130_as_sc_hs__inv_2 _3180_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\RAM[58][0] ),
    .Y(_1176_));
 sky130_as_sc_hs__nand4_2 _3181_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1175_),
    .B(\RAM[58][1] ),
    .C(_1176_),
    .Y(_1177_),
    .D(net8));
 sky130_as_sc_hs__inv_2 _3182_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\RAM[58][4] ),
    .Y(_1178_));
 sky130_as_sc_hs__nand3_2 _3183_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\RAM[58][5] ),
    .B(_1178_),
    .C(\RAM[58][3] ),
    .Y(_1179_));
 sky130_as_sc_hs__nor2_2 _3184_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1177_),
    .B(_1179_),
    .Y(HCF));
 sky130_as_sc_hs__buff_8 _3185_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1157_),
    .Y(_1180_));
 sky130_as_sc_hs__inv_2 _3186_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\ROM_spi_dat_out[0] ),
    .Y(_1181_));
 sky130_as_sc_hs__buff_4 _3187_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1123_),
    .Y(_1182_));
 sky130_as_sc_hs__inv_2 _3188_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\ROM_dest[0] ),
    .Y(_1183_));
 sky130_as_sc_hs__or2_2 _3189_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1183_),
    .B(_0669_),
    .Y(_1184_));
 sky130_as_sc_hs__clkbuff_4 _3190_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1184_),
    .Y(_1185_));
 sky130_as_sc_hs__mux2_2 _3191_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1185_),
    .B(_1182_),
    .A(_1181_),
    .Y(_1186_));
 sky130_as_sc_hs__nor2_2 _3192_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1180_),
    .B(_1186_),
    .Y(_0012_));
 sky130_as_sc_hs__inv_2 _3193_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\ROM_spi_dat_out[1] ),
    .Y(_1187_));
 sky130_as_sc_hs__mux2_2 _3194_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1185_),
    .B(_1129_),
    .A(_1187_),
    .Y(_1188_));
 sky130_as_sc_hs__nor2_2 _3195_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1180_),
    .B(_1188_),
    .Y(_0013_));
 sky130_as_sc_hs__mux2_2 _3196_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1185_),
    .B(net39),
    .A(\ROM_spi_dat_out[2] ),
    .Y(_1189_));
 sky130_as_sc_hs__and2_2 _3197_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net157),
    .B(_1189_),
    .Y(_1190_));
 sky130_as_sc_hs__buff_2 _3198_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1190_),
    .Y(_0014_));
 sky130_as_sc_hs__mux2_2 _3199_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1185_),
    .B(net35),
    .A(\ROM_spi_dat_out[3] ),
    .Y(_1191_));
 sky130_as_sc_hs__and2_2 _3200_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net157),
    .B(_1191_),
    .Y(_1192_));
 sky130_as_sc_hs__buff_2 _3201_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1192_),
    .Y(_0015_));
 sky130_as_sc_hs__mux2_2 _3202_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1185_),
    .B(net31),
    .A(\ROM_spi_dat_out[4] ),
    .Y(_1193_));
 sky130_as_sc_hs__and2_2 _3203_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net157),
    .B(_1193_),
    .Y(_1194_));
 sky130_as_sc_hs__buff_2 _3204_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1194_),
    .Y(_0016_));
 sky130_as_sc_hs__mux2_2 _3205_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1185_),
    .B(net29),
    .A(\ROM_spi_dat_out[5] ),
    .Y(_1195_));
 sky130_as_sc_hs__and2_2 _3206_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net157),
    .B(_1195_),
    .Y(_1196_));
 sky130_as_sc_hs__buff_2 _3207_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1196_),
    .Y(_0017_));
 sky130_as_sc_hs__mux2_2 _3208_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0653_),
    .B(net122),
    .A(_0999_),
    .Y(_1197_));
 sky130_as_sc_hs__mux2_2 _3209_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0660_),
    .B(\last_MAR[0] ),
    .A(net122),
    .Y(_1198_));
 sky130_as_sc_hs__ao22_2 _3210_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0926_),
    .C(_1198_),
    .B(_1197_),
    .D(_0657_),
    .Y(_1199_));
 sky130_as_sc_hs__ao22_2 _3211_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net123),
    .C(_1199_),
    .B(_1091_),
    .D(_1008_),
    .Y(_1200_));
 sky130_as_sc_hs__mux2_2 _3212_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0672_),
    .B(_1200_),
    .A(\ROM_spi_dat_out[0] ),
    .Y(_1201_));
 sky130_as_sc_hs__and2_2 _3213_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net151),
    .B(_1201_),
    .Y(_1202_));
 sky130_as_sc_hs__buff_2 _3214_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1202_),
    .Y(_0000_));
 sky130_as_sc_hs__mux2_2 _3215_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0653_),
    .B(net102),
    .A(_1084_),
    .Y(_1203_));
 sky130_as_sc_hs__mux2_2 _3216_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0660_),
    .B(\last_MAR[1] ),
    .A(net102),
    .Y(_1204_));
 sky130_as_sc_hs__ao22_2 _3217_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0534_),
    .C(_1204_),
    .B(_1203_),
    .D(_0657_),
    .Y(_1205_));
 sky130_as_sc_hs__ao22_2 _3218_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net102),
    .C(_1205_),
    .B(_1091_),
    .D(_0533_),
    .Y(_1206_));
 sky130_as_sc_hs__mux2_2 _3219_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0672_),
    .B(_1206_),
    .A(\ROM_spi_dat_out[1] ),
    .Y(_1207_));
 sky130_as_sc_hs__and2_2 _3220_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net151),
    .B(_1207_),
    .Y(_1208_));
 sky130_as_sc_hs__buff_2 _3221_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1208_),
    .Y(_0001_));
 sky130_as_sc_hs__nand2_2 _3222_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\instr_cycle[1] ),
    .B(_0655_),
    .Y(_1209_));
 sky130_as_sc_hs__or2_2 _3223_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net31),
    .B(net36),
    .Y(_1210_));
 sky130_as_sc_hs__nand2_4 _3224_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1150_),
    .B(net41),
    .Y(_1211_));
 sky130_as_sc_hs__or2_2 _3225_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1210_),
    .B(_1211_),
    .Y(_1212_));
 sky130_as_sc_hs__nor3_2 _3226_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0664_),
    .B(_1209_),
    .C(_1212_),
    .Y(_1213_));
 sky130_as_sc_hs__and2_2 _3227_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net148),
    .B(net21),
    .Y(_1214_));
 sky130_as_sc_hs__clkbuff_4 _3228_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1214_),
    .Y(_1215_));
 sky130_as_sc_hs__mux2_2 _3229_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net48),
    .B(net132),
    .A(\B[0] ),
    .Y(_1216_));
 sky130_as_sc_hs__and2_2 _3230_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1215_),
    .B(_1216_),
    .Y(_1217_));
 sky130_as_sc_hs__buff_2 _3231_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1217_),
    .Y(_1218_));
 sky130_as_sc_hs__buff_4 _3232_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1218_),
    .Y(_1219_));
 sky130_as_sc_hs__nand2_2 _3233_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net148),
    .B(net21),
    .Y(_1220_));
 sky130_as_sc_hs__or2_2 _3234_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net88),
    .B(_1220_),
    .Y(_1221_));
 sky130_as_sc_hs__or2_2 _3235_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0627_),
    .B(_1221_),
    .Y(_1222_));
 sky130_as_sc_hs__clkbuff_11 _3236_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1222_),
    .Y(_1223_));
 sky130_as_sc_hs__nand2_2 _3237_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0632_),
    .B(_1214_),
    .Y(_1224_));
 sky130_as_sc_hs__buff_6 _3238_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1224_),
    .Y(_1225_));
 sky130_as_sc_hs__nor2_4 _3239_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1223_),
    .B(_1225_),
    .Y(_1226_));
 sky130_as_sc_hs__mux2_2 _3240_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1226_),
    .B(_1219_),
    .A(net304),
    .Y(_1227_));
 sky130_as_sc_hs__buff_2 _3241_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1227_),
    .Y(_0024_));
 sky130_as_sc_hs__mux2_2 _3242_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net48),
    .B(net131),
    .A(\B[1] ),
    .Y(_1228_));
 sky130_as_sc_hs__and2_2 _3243_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1215_),
    .B(_1228_),
    .Y(_1229_));
 sky130_as_sc_hs__buff_2 _3244_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1229_),
    .Y(_1230_));
 sky130_as_sc_hs__buff_2 _3245_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1230_),
    .Y(_1231_));
 sky130_as_sc_hs__mux2_2 _3246_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1226_),
    .B(_1231_),
    .A(net283),
    .Y(_1232_));
 sky130_as_sc_hs__buff_2 _3247_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1232_),
    .Y(_0025_));
 sky130_as_sc_hs__mux2_2 _3248_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net48),
    .B(net129),
    .A(\B[2] ),
    .Y(_1233_));
 sky130_as_sc_hs__and2_2 _3249_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1215_),
    .B(_1233_),
    .Y(_1234_));
 sky130_as_sc_hs__buff_2 _3250_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1234_),
    .Y(_1235_));
 sky130_as_sc_hs__clkbuff_4 _3251_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1235_),
    .Y(_1236_));
 sky130_as_sc_hs__mux2_2 _3252_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1226_),
    .B(_1236_),
    .A(net322),
    .Y(_1237_));
 sky130_as_sc_hs__buff_2 _3253_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1237_),
    .Y(_0026_));
 sky130_as_sc_hs__mux2_2 _3254_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net48),
    .B(\A[3] ),
    .A(\B[3] ),
    .Y(_1238_));
 sky130_as_sc_hs__and2_2 _3255_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1215_),
    .B(_1238_),
    .Y(_1239_));
 sky130_as_sc_hs__clkbuff_4 _3256_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1239_),
    .Y(_1240_));
 sky130_as_sc_hs__clkbuff_4 _3257_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1240_),
    .Y(_1241_));
 sky130_as_sc_hs__mux2_2 _3258_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1226_),
    .B(_1241_),
    .A(net355),
    .Y(_1242_));
 sky130_as_sc_hs__buff_2 _3259_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1242_),
    .Y(_0027_));
 sky130_as_sc_hs__inv_2 _3260_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\B[4] ),
    .Y(_1243_));
 sky130_as_sc_hs__inv_2 _3261_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net126),
    .Y(_1244_));
 sky130_as_sc_hs__mux2_2 _3262_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net48),
    .B(_1244_),
    .A(_1243_),
    .Y(_1245_));
 sky130_as_sc_hs__nor2_4 _3263_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1220_),
    .B(_1245_),
    .Y(_1246_));
 sky130_as_sc_hs__buff_2 _3264_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1246_),
    .Y(_1247_));
 sky130_as_sc_hs__clkbuff_4 _3265_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1247_),
    .Y(_1248_));
 sky130_as_sc_hs__mux2_2 _3266_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1226_),
    .B(_1248_),
    .A(net578),
    .Y(_1249_));
 sky130_as_sc_hs__buff_2 _3267_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1249_),
    .Y(_0028_));
 sky130_as_sc_hs__mux2_2 _3268_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net48),
    .B(net124),
    .A(\B[5] ),
    .Y(_1250_));
 sky130_as_sc_hs__and2_2 _3269_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1214_),
    .B(_1250_),
    .Y(_1251_));
 sky130_as_sc_hs__buff_2 _3270_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1251_),
    .Y(_1252_));
 sky130_as_sc_hs__clkbuff_4 _3271_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1252_),
    .Y(_1253_));
 sky130_as_sc_hs__mux2_2 _3272_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1226_),
    .B(_1253_),
    .A(net553),
    .Y(_1254_));
 sky130_as_sc_hs__buff_2 _3273_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1254_),
    .Y(_0029_));
 sky130_as_sc_hs__or2_2 _3274_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1053_),
    .B(_1221_),
    .Y(_1255_));
 sky130_as_sc_hs__clkbuff_11 _3275_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1255_),
    .Y(_1256_));
 sky130_as_sc_hs__nor2_4 _3276_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1225_),
    .B(_1256_),
    .Y(_1257_));
 sky130_as_sc_hs__mux2_2 _3277_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1257_),
    .B(_1219_),
    .A(net293),
    .Y(_1258_));
 sky130_as_sc_hs__buff_2 _3278_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1258_),
    .Y(_0030_));
 sky130_as_sc_hs__mux2_2 _3279_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1257_),
    .B(_1231_),
    .A(net352),
    .Y(_1259_));
 sky130_as_sc_hs__buff_2 _3280_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1259_),
    .Y(_0031_));
 sky130_as_sc_hs__mux2_2 _3281_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1257_),
    .B(_1236_),
    .A(net505),
    .Y(_1260_));
 sky130_as_sc_hs__buff_2 _3282_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1260_),
    .Y(_0032_));
 sky130_as_sc_hs__mux2_2 _3283_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1257_),
    .B(_1241_),
    .A(net215),
    .Y(_1261_));
 sky130_as_sc_hs__buff_2 _3284_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1261_),
    .Y(_0033_));
 sky130_as_sc_hs__mux2_2 _3285_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1257_),
    .B(_1248_),
    .A(net427),
    .Y(_1262_));
 sky130_as_sc_hs__buff_2 _3286_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1262_),
    .Y(_0034_));
 sky130_as_sc_hs__mux2_2 _3287_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1257_),
    .B(_1253_),
    .A(net565),
    .Y(_1263_));
 sky130_as_sc_hs__buff_2 _3288_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1263_),
    .Y(_0035_));
 sky130_as_sc_hs__nand2_2 _3289_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net88),
    .B(_1214_),
    .Y(_1264_));
 sky130_as_sc_hs__or2_2 _3290_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0627_),
    .B(_1264_),
    .Y(_1265_));
 sky130_as_sc_hs__clkbuff_11 _3291_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1265_),
    .Y(_1266_));
 sky130_as_sc_hs__nor2_4 _3292_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0638_),
    .B(_1266_),
    .Y(_1267_));
 sky130_as_sc_hs__mux2_2 _3293_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1267_),
    .B(_1219_),
    .A(net229),
    .Y(_1268_));
 sky130_as_sc_hs__buff_2 _3294_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1268_),
    .Y(_0036_));
 sky130_as_sc_hs__mux2_2 _3295_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1267_),
    .B(_1231_),
    .A(net581),
    .Y(_1269_));
 sky130_as_sc_hs__buff_2 _3296_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1269_),
    .Y(_0037_));
 sky130_as_sc_hs__mux2_2 _3297_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1267_),
    .B(_1236_),
    .A(net587),
    .Y(_1270_));
 sky130_as_sc_hs__buff_2 _3298_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1270_),
    .Y(_0038_));
 sky130_as_sc_hs__mux2_2 _3299_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1267_),
    .B(_1241_),
    .A(net521),
    .Y(_1271_));
 sky130_as_sc_hs__buff_2 _3300_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1271_),
    .Y(_0039_));
 sky130_as_sc_hs__mux2_2 _3301_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1267_),
    .B(_1248_),
    .A(net580),
    .Y(_1272_));
 sky130_as_sc_hs__buff_2 _3302_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1272_),
    .Y(_0040_));
 sky130_as_sc_hs__mux2_2 _3303_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1267_),
    .B(_1253_),
    .A(net573),
    .Y(_1273_));
 sky130_as_sc_hs__buff_2 _3304_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1273_),
    .Y(_0041_));
 sky130_as_sc_hs__or2_4 _3305_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1056_),
    .B(_1221_),
    .Y(_1274_));
 sky130_as_sc_hs__buff_11 _3306_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1274_),
    .Y(_1275_));
 sky130_as_sc_hs__nand2_4 _3307_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0610_),
    .B(_1215_),
    .Y(_1276_));
 sky130_as_sc_hs__nor2_4 _3308_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1275_),
    .B(_1276_),
    .Y(_1277_));
 sky130_as_sc_hs__mux2_2 _3309_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1277_),
    .B(_1219_),
    .A(net198),
    .Y(_1278_));
 sky130_as_sc_hs__buff_2 _3310_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1278_),
    .Y(_0042_));
 sky130_as_sc_hs__mux2_2 _3311_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1277_),
    .B(_1231_),
    .A(net363),
    .Y(_1279_));
 sky130_as_sc_hs__buff_2 _3312_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1279_),
    .Y(_0043_));
 sky130_as_sc_hs__mux2_2 _3313_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1277_),
    .B(_1236_),
    .A(net326),
    .Y(_1280_));
 sky130_as_sc_hs__buff_2 _3314_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1280_),
    .Y(_0044_));
 sky130_as_sc_hs__mux2_2 _3315_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1277_),
    .B(_1241_),
    .A(net468),
    .Y(_1281_));
 sky130_as_sc_hs__buff_2 _3316_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1281_),
    .Y(_0045_));
 sky130_as_sc_hs__mux2_2 _3317_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1277_),
    .B(_1248_),
    .A(net436),
    .Y(_1282_));
 sky130_as_sc_hs__buff_2 _3318_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1282_),
    .Y(_0046_));
 sky130_as_sc_hs__mux2_2 _3319_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1277_),
    .B(_1253_),
    .A(net525),
    .Y(_1283_));
 sky130_as_sc_hs__buff_2 _3320_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1283_),
    .Y(_0047_));
 sky130_as_sc_hs__inv_2 _3321_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net145),
    .Y(_1284_));
 sky130_as_sc_hs__buff_2 _3322_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0668_),
    .Y(_1285_));
 sky130_as_sc_hs__nor2_2 _3323_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1138_),
    .B(_1123_),
    .Y(_1286_));
 sky130_as_sc_hs__ao21_2 _3324_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1162_),
    .B(_1286_),
    .C(_1169_),
    .Y(_1287_));
 sky130_as_sc_hs__ao21_2 _3325_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1139_),
    .B(_1152_),
    .C(net28),
    .Y(_1288_));
 sky130_as_sc_hs__nand2_2 _3326_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1151_),
    .B(_1288_),
    .Y(_1289_));
 sky130_as_sc_hs__ao31_4 _3327_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1161_),
    .B(_1287_),
    .C(_1289_),
    .D(net139),
    .Y(_1290_));
 sky130_as_sc_hs__or2_2 _3328_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0531_),
    .B(_1290_),
    .Y(_1291_));
 sky130_as_sc_hs__buff_2 _3329_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0530_),
    .Y(_1292_));
 sky130_as_sc_hs__clkbuff_4 _3330_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1292_),
    .Y(_1293_));
 sky130_as_sc_hs__ao21_2 _3331_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net145),
    .B(_1293_),
    .C(_1156_),
    .Y(_1294_));
 sky130_as_sc_hs__ao31_2 _3332_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1284_),
    .B(_1285_),
    .C(_1291_),
    .D(_1294_),
    .Y(_1295_));
 sky130_as_sc_hs__buff_2 _3333_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1295_),
    .Y(_0048_));
 sky130_as_sc_hs__inv_2 _3334_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\mem_cycle[1] ),
    .Y(_1296_));
 sky130_as_sc_hs__nand2_2 _3335_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net144),
    .B(_0668_),
    .Y(_1297_));
 sky130_as_sc_hs__xnor2_2 _3336_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1296_),
    .Y(_1298_),
    .B(_1297_));
 sky130_as_sc_hs__nor2_2 _3337_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1180_),
    .B(_1298_),
    .Y(_0049_));
 sky130_as_sc_hs__xnor2_2 _3338_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_addr[10] ),
    .Y(_1299_),
    .B(\ROM_addr_buff[10] ));
 sky130_as_sc_hs__nand4_2 _3339_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_addr[3] ),
    .B(\last_addr[2] ),
    .C(\last_addr[1] ),
    .Y(_1300_),
    .D(\last_addr[0] ));
 sky130_as_sc_hs__nand2_2 _3340_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_addr[5] ),
    .B(\last_addr[4] ),
    .Y(_1301_));
 sky130_as_sc_hs__or2_2 _3341_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1300_),
    .B(_1301_),
    .Y(_1302_));
 sky130_as_sc_hs__nand2_2 _3342_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_addr[7] ),
    .B(\last_addr[6] ),
    .Y(_1303_));
 sky130_as_sc_hs__nor2_2 _3343_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1302_),
    .B(_1303_),
    .Y(_1304_));
 sky130_as_sc_hs__nand2_2 _3344_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_addr[8] ),
    .B(_1304_),
    .Y(_1305_));
 sky130_as_sc_hs__inv_2 _3345_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\ROM_addr_buff[11] ),
    .Y(_1306_));
 sky130_as_sc_hs__nor2_2 _3346_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_addr[11] ),
    .B(_1306_),
    .Y(_1307_));
 sky130_as_sc_hs__oai21_2 _3347_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1305_),
    .B(_1307_),
    .C(net27),
    .Y(_1308_));
 sky130_as_sc_hs__and2_2 _3348_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1299_),
    .B(_1308_),
    .Y(_1309_));
 sky130_as_sc_hs__oa21_2 _3349_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_addr[11] ),
    .B(_1306_),
    .C(_1299_),
    .Y(_1310_));
 sky130_as_sc_hs__nor3_2 _3350_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net27),
    .B(_1305_),
    .C(_1299_),
    .Y(_1311_));
 sky130_as_sc_hs__ao31_2 _3351_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net27),
    .B(_1305_),
    .C(_1310_),
    .D(_1311_),
    .Y(_1312_));
 sky130_as_sc_hs__mux2_2 _3352_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(\last_addr[9] ),
    .B(_1312_),
    .A(_1309_),
    .Y(_1313_));
 sky130_as_sc_hs__xnor2_2 _3353_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_addr[7] ),
    .Y(_1314_),
    .B(\ROM_addr_buff[7] ));
 sky130_as_sc_hs__nand2b_2 _3354_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(\last_addr[6] ),
    .Y(_1315_),
    .A(\ROM_addr_buff[6] ));
 sky130_as_sc_hs__nand2b_2 _3355_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(\ROM_addr_buff[6] ),
    .Y(_1316_),
    .A(\last_addr[6] ));
 sky130_as_sc_hs__and2_2 _3356_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1315_),
    .B(_1316_),
    .Y(_1317_));
 sky130_as_sc_hs__mux2_2 _3357_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1314_),
    .B(_1316_),
    .A(_1315_),
    .Y(_1318_));
 sky130_as_sc_hs__nor2_2 _3358_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1302_),
    .B(_1318_),
    .Y(_1319_));
 sky130_as_sc_hs__ao31_2 _3359_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1302_),
    .B(_1314_),
    .C(_1317_),
    .D(_1319_),
    .Y(_1320_));
 sky130_as_sc_hs__xnor2_2 _3360_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_addr_buff[8] ),
    .Y(_1321_),
    .B(_1304_));
 sky130_as_sc_hs__nor2_2 _3361_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_addr[9] ),
    .B(\ROM_addr_buff[9] ),
    .Y(_1322_));
 sky130_as_sc_hs__ao31_2 _3362_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_addr[11] ),
    .B(\last_addr[10] ),
    .C(\last_addr[9] ),
    .D(_1322_),
    .Y(_1323_));
 sky130_as_sc_hs__nor2_2 _3363_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\ROM_addr_buff[8] ),
    .B(_1323_),
    .Y(_1324_));
 sky130_as_sc_hs__mux2_2 _3364_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1304_),
    .B(_1324_),
    .A(\ROM_addr_buff[8] ),
    .Y(_1325_));
 sky130_as_sc_hs__mux2_2 _3365_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(\last_addr[8] ),
    .B(_1325_),
    .A(_1321_),
    .Y(_1326_));
 sky130_as_sc_hs__inv_2 _3366_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\last_addr[4] ),
    .Y(_1327_));
 sky130_as_sc_hs__xnor2_2 _3367_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_addr[5] ),
    .Y(_1328_),
    .B(\ROM_addr_buff[5] ));
 sky130_as_sc_hs__nor3_2 _3368_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1327_),
    .B(\ROM_addr_buff[4] ),
    .C(_1328_),
    .Y(_1329_));
 sky130_as_sc_hs__nand3_2 _3369_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1327_),
    .B(\ROM_addr_buff[4] ),
    .C(_1328_),
    .Y(_1330_));
 sky130_as_sc_hs__ao21b_2 _3370_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1329_),
    .B(_1330_),
    .C(_1300_),
    .Y(_1331_));
 sky130_as_sc_hs__xnor2_2 _3371_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_addr[4] ),
    .Y(_1332_),
    .B(\ROM_addr_buff[4] ));
 sky130_as_sc_hs__nand3_2 _3372_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1300_),
    .B(_1328_),
    .C(_1332_),
    .Y(_1333_));
 sky130_as_sc_hs__nand2_2 _3373_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_addr[10] ),
    .B(\last_addr[9] ),
    .Y(_1334_));
 sky130_as_sc_hs__nor2_2 _3374_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net27),
    .B(_1334_),
    .Y(_1335_));
 sky130_as_sc_hs__nor2_2 _3375_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_addr[11] ),
    .B(_1335_),
    .Y(_1336_));
 sky130_as_sc_hs__inv_2 _3376_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\last_addr[2] ),
    .Y(_1337_));
 sky130_as_sc_hs__nor2_2 _3377_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1337_),
    .B(\ROM_addr_buff[2] ),
    .Y(_1338_));
 sky130_as_sc_hs__nand2_2 _3378_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_addr[1] ),
    .B(\last_addr[0] ),
    .Y(_1339_));
 sky130_as_sc_hs__ao21_2 _3379_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1337_),
    .B(\ROM_addr_buff[2] ),
    .C(_1339_),
    .Y(_1340_));
 sky130_as_sc_hs__xnor2_2 _3380_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_addr[3] ),
    .Y(_1341_),
    .B(\ROM_addr_buff[3] ));
 sky130_as_sc_hs__mux2_2 _3381_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1341_),
    .B(_1340_),
    .A(_1338_),
    .Y(_1342_));
 sky130_as_sc_hs__aoi211_2 _3382_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1334_),
    .C(_1284_),
    .D(_0531_),
    .Y(_1343_),
    .A(_1307_));
 sky130_as_sc_hs__iao211_2 _3383_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_addr_buff[11] ),
    .B(_1336_),
    .C(_1342_),
    .D(_1343_),
    .Y(_1344_));
 sky130_as_sc_hs__xnor2_2 _3384_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_addr[2] ),
    .Y(_1345_),
    .B(\ROM_addr_buff[2] ));
 sky130_as_sc_hs__inv_2 _3385_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\last_addr[0] ),
    .Y(_1346_));
 sky130_as_sc_hs__xnor2_2 _3386_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_addr[1] ),
    .Y(_1347_),
    .B(\ROM_addr_buff[1] ));
 sky130_as_sc_hs__nand2b_2 _3387_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .B(\ROM_addr_buff[1] ),
    .Y(_1348_),
    .A(\last_addr[1] ));
 sky130_as_sc_hs__nor3_2 _3388_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1346_),
    .B(\ROM_addr_buff[0] ),
    .C(_1348_),
    .Y(_1349_));
 sky130_as_sc_hs__ao31_2 _3389_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1346_),
    .B(\ROM_addr_buff[0] ),
    .C(_1347_),
    .D(_1349_),
    .Y(_1350_));
 sky130_as_sc_hs__nor3_2 _3390_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\ROM_addr_buff[1] ),
    .B(\ROM_addr_buff[0] ),
    .C(_1339_),
    .Y(_1351_));
 sky130_as_sc_hs__aoi21_2 _3391_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1345_),
    .B(_1350_),
    .C(_1351_),
    .Y(_1352_));
 sky130_as_sc_hs__aoi211_2 _3392_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1333_),
    .C(_1344_),
    .D(_1352_),
    .Y(_1353_),
    .A(_1331_));
 sky130_as_sc_hs__nand4_2 _3393_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1313_),
    .B(_1320_),
    .C(_1326_),
    .Y(_1354_),
    .D(_1353_));
 sky130_as_sc_hs__oa21_2 _3394_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1296_),
    .B(_1284_),
    .C(_1354_),
    .Y(_1355_));
 sky130_as_sc_hs__aoi211_2 _3395_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1284_),
    .C(_1293_),
    .D(_1355_),
    .Y(_1356_),
    .A(_1296_));
 sky130_as_sc_hs__iao211_2 _3396_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net143),
    .B(_1356_),
    .C(_0669_),
    .D(net152),
    .Y(_1357_));
 sky130_as_sc_hs__inv_2 _3397_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_1357_),
    .Y(_0050_));
 sky130_as_sc_hs__nor2_4 _3398_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1225_),
    .B(_1266_),
    .Y(_1358_));
 sky130_as_sc_hs__mux2_2 _3399_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1358_),
    .B(_1219_),
    .A(net424),
    .Y(_1359_));
 sky130_as_sc_hs__buff_2 _3400_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1359_),
    .Y(_0051_));
 sky130_as_sc_hs__mux2_2 _3401_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1358_),
    .B(_1231_),
    .A(net277),
    .Y(_1360_));
 sky130_as_sc_hs__buff_2 _3402_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1360_),
    .Y(_0052_));
 sky130_as_sc_hs__mux2_2 _3403_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1358_),
    .B(_1236_),
    .A(net332),
    .Y(_1361_));
 sky130_as_sc_hs__buff_2 _3404_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1361_),
    .Y(_0053_));
 sky130_as_sc_hs__mux2_2 _3405_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1358_),
    .B(_1241_),
    .A(net540),
    .Y(_1362_));
 sky130_as_sc_hs__buff_2 _3406_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1362_),
    .Y(_0054_));
 sky130_as_sc_hs__mux2_2 _3407_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1358_),
    .B(_1248_),
    .A(net354),
    .Y(_1363_));
 sky130_as_sc_hs__buff_2 _3408_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1363_),
    .Y(_0055_));
 sky130_as_sc_hs__mux2_2 _3409_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1358_),
    .B(_1253_),
    .A(net547),
    .Y(_1364_));
 sky130_as_sc_hs__buff_2 _3410_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1364_),
    .Y(_0056_));
 sky130_as_sc_hs__or2_2 _3411_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1056_),
    .B(_1264_),
    .Y(_1365_));
 sky130_as_sc_hs__clkbuff_11 _3412_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1365_),
    .Y(_1366_));
 sky130_as_sc_hs__nand2_2 _3413_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0588_),
    .B(_1214_),
    .Y(_1367_));
 sky130_as_sc_hs__or2_2 _3414_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0609_),
    .B(_1367_),
    .Y(_1368_));
 sky130_as_sc_hs__buff_6 _3415_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1368_),
    .Y(_1369_));
 sky130_as_sc_hs__nor2_4 _3416_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1366_),
    .B(_1369_),
    .Y(_1370_));
 sky130_as_sc_hs__mux2_2 _3417_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1370_),
    .B(_1219_),
    .A(net451),
    .Y(_1371_));
 sky130_as_sc_hs__buff_2 _3418_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1371_),
    .Y(_0057_));
 sky130_as_sc_hs__mux2_2 _3419_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1370_),
    .B(_1231_),
    .A(net294),
    .Y(_1372_));
 sky130_as_sc_hs__buff_2 _3420_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1372_),
    .Y(_0058_));
 sky130_as_sc_hs__mux2_2 _3421_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1370_),
    .B(_1236_),
    .A(net506),
    .Y(_1373_));
 sky130_as_sc_hs__buff_2 _3422_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1373_),
    .Y(_0059_));
 sky130_as_sc_hs__mux2_2 _3423_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1370_),
    .B(_1241_),
    .A(net317),
    .Y(_1374_));
 sky130_as_sc_hs__buff_2 _3424_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1374_),
    .Y(_0060_));
 sky130_as_sc_hs__mux2_2 _3425_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1370_),
    .B(_1248_),
    .A(net585),
    .Y(_1375_));
 sky130_as_sc_hs__buff_2 _3426_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1375_),
    .Y(_0061_));
 sky130_as_sc_hs__mux2_2 _3427_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1370_),
    .B(_1253_),
    .A(net426),
    .Y(_1376_));
 sky130_as_sc_hs__buff_2 _3428_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1376_),
    .Y(_0062_));
 sky130_as_sc_hs__and2_4 _3429_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0639_),
    .B(_1215_),
    .Y(_1377_));
 sky130_as_sc_hs__nor2_4 _3430_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1225_),
    .B(_1377_),
    .Y(_1378_));
 sky130_as_sc_hs__mux2_2 _3431_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1378_),
    .B(_1219_),
    .A(net362),
    .Y(_1379_));
 sky130_as_sc_hs__buff_2 _3432_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1379_),
    .Y(_0063_));
 sky130_as_sc_hs__mux2_2 _3433_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1378_),
    .B(_1231_),
    .A(net419),
    .Y(_1380_));
 sky130_as_sc_hs__buff_2 _3434_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1380_),
    .Y(_0064_));
 sky130_as_sc_hs__mux2_2 _3435_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1378_),
    .B(_1236_),
    .A(net325),
    .Y(_1381_));
 sky130_as_sc_hs__buff_2 _3436_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1381_),
    .Y(_0065_));
 sky130_as_sc_hs__mux2_2 _3437_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1378_),
    .B(_1241_),
    .A(net487),
    .Y(_1382_));
 sky130_as_sc_hs__buff_2 _3438_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1382_),
    .Y(_0066_));
 sky130_as_sc_hs__mux2_2 _3439_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1378_),
    .B(_1248_),
    .A(net455),
    .Y(_1383_));
 sky130_as_sc_hs__buff_2 _3440_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1383_),
    .Y(_0067_));
 sky130_as_sc_hs__mux2_2 _3441_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1378_),
    .B(_1253_),
    .A(net498),
    .Y(_1384_));
 sky130_as_sc_hs__buff_2 _3442_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1384_),
    .Y(_0068_));
 sky130_as_sc_hs__buff_4 _3443_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1218_),
    .Y(_1385_));
 sky130_as_sc_hs__or2_2 _3444_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0606_),
    .B(_1367_),
    .Y(_1386_));
 sky130_as_sc_hs__buff_6 _3445_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1386_),
    .Y(_1387_));
 sky130_as_sc_hs__nor2_4 _3446_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1256_),
    .B(_1387_),
    .Y(_1388_));
 sky130_as_sc_hs__mux2_2 _3447_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1388_),
    .B(_1385_),
    .A(net527),
    .Y(_1389_));
 sky130_as_sc_hs__buff_2 _3448_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1389_),
    .Y(_0069_));
 sky130_as_sc_hs__clkbuff_4 _3449_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1230_),
    .Y(_1390_));
 sky130_as_sc_hs__mux2_2 _3450_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1388_),
    .B(_1390_),
    .A(net366),
    .Y(_1391_));
 sky130_as_sc_hs__buff_2 _3451_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1391_),
    .Y(_0070_));
 sky130_as_sc_hs__clkbuff_4 _3452_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1235_),
    .Y(_1392_));
 sky130_as_sc_hs__mux2_2 _3453_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1388_),
    .B(_1392_),
    .A(net481),
    .Y(_1393_));
 sky130_as_sc_hs__buff_2 _3454_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1393_),
    .Y(_0071_));
 sky130_as_sc_hs__buff_4 _3455_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1240_),
    .Y(_1394_));
 sky130_as_sc_hs__mux2_2 _3456_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1388_),
    .B(_1394_),
    .A(net558),
    .Y(_1395_));
 sky130_as_sc_hs__buff_2 _3457_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1395_),
    .Y(_0072_));
 sky130_as_sc_hs__buff_4 _3458_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1247_),
    .Y(_1396_));
 sky130_as_sc_hs__mux2_2 _3459_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1388_),
    .B(_1396_),
    .A(net471),
    .Y(_1397_));
 sky130_as_sc_hs__buff_2 _3460_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1397_),
    .Y(_0073_));
 sky130_as_sc_hs__buff_4 _3461_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1252_),
    .Y(_1398_));
 sky130_as_sc_hs__mux2_2 _3462_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1388_),
    .B(_1398_),
    .A(net397),
    .Y(_1399_));
 sky130_as_sc_hs__buff_2 _3463_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1399_),
    .Y(_0074_));
 sky130_as_sc_hs__nand2_4 _3464_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net141),
    .B(_0989_),
    .Y(_1400_));
 sky130_as_sc_hs__or2_2 _3465_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0625_),
    .B(_1221_),
    .Y(_1401_));
 sky130_as_sc_hs__clkbuff_11 _3466_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1401_),
    .Y(_1402_));
 sky130_as_sc_hs__nor2_4 _3467_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1400_),
    .B(_1402_),
    .Y(_1403_));
 sky130_as_sc_hs__mux2_2 _3468_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1403_),
    .B(_1385_),
    .A(net241),
    .Y(_1404_));
 sky130_as_sc_hs__buff_2 _3469_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1404_),
    .Y(_0075_));
 sky130_as_sc_hs__mux2_2 _3470_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1403_),
    .B(_1390_),
    .A(net311),
    .Y(_1405_));
 sky130_as_sc_hs__buff_2 _3471_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1405_),
    .Y(_0076_));
 sky130_as_sc_hs__mux2_2 _3472_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1403_),
    .B(_1392_),
    .A(net287),
    .Y(_1406_));
 sky130_as_sc_hs__buff_2 _3473_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1406_),
    .Y(_0077_));
 sky130_as_sc_hs__mux2_2 _3474_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1403_),
    .B(_1394_),
    .A(net369),
    .Y(_1407_));
 sky130_as_sc_hs__buff_2 _3475_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1407_),
    .Y(_0078_));
 sky130_as_sc_hs__mux2_2 _3476_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1403_),
    .B(_1396_),
    .A(net526),
    .Y(_1408_));
 sky130_as_sc_hs__buff_2 _3477_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1408_),
    .Y(_0079_));
 sky130_as_sc_hs__mux2_2 _3478_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1403_),
    .B(_1398_),
    .A(net379),
    .Y(_1409_));
 sky130_as_sc_hs__buff_2 _3479_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1409_),
    .Y(_0080_));
 sky130_as_sc_hs__nand2_2 _3480_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0590_),
    .B(_1215_),
    .Y(_1410_));
 sky130_as_sc_hs__buff_6 _3481_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1410_),
    .Y(_1411_));
 sky130_as_sc_hs__nor2_4 _3482_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1377_),
    .B(_1411_),
    .Y(_1412_));
 sky130_as_sc_hs__mux2_2 _3483_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1412_),
    .B(_1385_),
    .A(net246),
    .Y(_1413_));
 sky130_as_sc_hs__buff_2 _3484_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1413_),
    .Y(_0081_));
 sky130_as_sc_hs__mux2_2 _3485_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1412_),
    .B(_1390_),
    .A(net351),
    .Y(_1414_));
 sky130_as_sc_hs__buff_2 _3486_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1414_),
    .Y(_0082_));
 sky130_as_sc_hs__mux2_2 _3487_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1412_),
    .B(_1392_),
    .A(net422),
    .Y(_1415_));
 sky130_as_sc_hs__buff_2 _3488_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1415_),
    .Y(_0083_));
 sky130_as_sc_hs__mux2_2 _3489_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1412_),
    .B(_1394_),
    .A(net516),
    .Y(_1416_));
 sky130_as_sc_hs__buff_2 _3490_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1416_),
    .Y(_0084_));
 sky130_as_sc_hs__mux2_2 _3491_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1412_),
    .B(_1396_),
    .A(net353),
    .Y(_1417_));
 sky130_as_sc_hs__buff_2 _3492_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1417_),
    .Y(_0085_));
 sky130_as_sc_hs__mux2_2 _3493_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1412_),
    .B(_1398_),
    .A(net296),
    .Y(_1418_));
 sky130_as_sc_hs__buff_2 _3494_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1418_),
    .Y(_0086_));
 sky130_as_sc_hs__nor2_4 _3495_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0607_),
    .B(_1220_),
    .Y(_1419_));
 sky130_as_sc_hs__nor2_4 _3496_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1275_),
    .B(_1419_),
    .Y(_1420_));
 sky130_as_sc_hs__mux2_2 _3497_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1420_),
    .B(_1385_),
    .A(net192),
    .Y(_1421_));
 sky130_as_sc_hs__buff_2 _3498_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1421_),
    .Y(_0087_));
 sky130_as_sc_hs__mux2_2 _3499_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1420_),
    .B(_1390_),
    .A(net259),
    .Y(_1422_));
 sky130_as_sc_hs__buff_2 _3500_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1422_),
    .Y(_0088_));
 sky130_as_sc_hs__mux2_2 _3501_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1420_),
    .B(_1392_),
    .A(net404),
    .Y(_1423_));
 sky130_as_sc_hs__buff_2 _3502_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1423_),
    .Y(_0089_));
 sky130_as_sc_hs__mux2_2 _3503_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1420_),
    .B(_1394_),
    .A(net358),
    .Y(_1424_));
 sky130_as_sc_hs__buff_2 _3504_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1424_),
    .Y(_0090_));
 sky130_as_sc_hs__mux2_2 _3505_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1420_),
    .B(_1396_),
    .A(net195),
    .Y(_1425_));
 sky130_as_sc_hs__buff_2 _3506_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1425_),
    .Y(_0091_));
 sky130_as_sc_hs__mux2_2 _3507_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1420_),
    .B(_1398_),
    .A(net203),
    .Y(_1426_));
 sky130_as_sc_hs__buff_2 _3508_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1426_),
    .Y(_0092_));
 sky130_as_sc_hs__or2_2 _3509_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0589_),
    .B(_1367_),
    .Y(_1427_));
 sky130_as_sc_hs__buff_6 _3510_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1427_),
    .Y(_1428_));
 sky130_as_sc_hs__nor2_4 _3511_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1223_),
    .B(_1428_),
    .Y(_1429_));
 sky130_as_sc_hs__mux2_2 _3512_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1429_),
    .B(_1385_),
    .A(net227),
    .Y(_1430_));
 sky130_as_sc_hs__buff_2 _3513_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1430_),
    .Y(_0093_));
 sky130_as_sc_hs__mux2_2 _3514_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1429_),
    .B(_1390_),
    .A(net344),
    .Y(_1431_));
 sky130_as_sc_hs__buff_2 _3515_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1431_),
    .Y(_0094_));
 sky130_as_sc_hs__mux2_2 _3516_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1429_),
    .B(_1392_),
    .A(net459),
    .Y(_1432_));
 sky130_as_sc_hs__buff_2 _3517_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1432_),
    .Y(_0095_));
 sky130_as_sc_hs__mux2_2 _3518_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1429_),
    .B(_1394_),
    .A(net338),
    .Y(_1433_));
 sky130_as_sc_hs__buff_2 _3519_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1433_),
    .Y(_0096_));
 sky130_as_sc_hs__mux2_2 _3520_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1429_),
    .B(_1396_),
    .A(net458),
    .Y(_1434_));
 sky130_as_sc_hs__buff_2 _3521_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1434_),
    .Y(_0097_));
 sky130_as_sc_hs__mux2_2 _3522_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1429_),
    .B(_1398_),
    .A(net290),
    .Y(_1435_));
 sky130_as_sc_hs__buff_2 _3523_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1435_),
    .Y(_0098_));
 sky130_as_sc_hs__nor2_4 _3524_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1400_),
    .B(_1266_),
    .Y(_1436_));
 sky130_as_sc_hs__mux2_2 _3525_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1436_),
    .B(_1385_),
    .A(net328),
    .Y(_1437_));
 sky130_as_sc_hs__buff_2 _3526_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1437_),
    .Y(_0099_));
 sky130_as_sc_hs__mux2_2 _3527_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1436_),
    .B(_1390_),
    .A(net257),
    .Y(_1438_));
 sky130_as_sc_hs__buff_2 _3528_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1438_),
    .Y(_0100_));
 sky130_as_sc_hs__mux2_2 _3529_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1436_),
    .B(_1392_),
    .A(net269),
    .Y(_1439_));
 sky130_as_sc_hs__buff_2 _3530_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1439_),
    .Y(_0101_));
 sky130_as_sc_hs__mux2_2 _3531_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1436_),
    .B(_1394_),
    .A(net224),
    .Y(_1440_));
 sky130_as_sc_hs__buff_2 _3532_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1440_),
    .Y(_0102_));
 sky130_as_sc_hs__mux2_2 _3533_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1436_),
    .B(_1396_),
    .A(net515),
    .Y(_1441_));
 sky130_as_sc_hs__buff_2 _3534_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1441_),
    .Y(_0103_));
 sky130_as_sc_hs__mux2_2 _3535_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1436_),
    .B(_1398_),
    .A(net394),
    .Y(_1442_));
 sky130_as_sc_hs__buff_2 _3536_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1442_),
    .Y(_0104_));
 sky130_as_sc_hs__nor2_4 _3537_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1276_),
    .B(_1377_),
    .Y(_1443_));
 sky130_as_sc_hs__mux2_2 _3538_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1443_),
    .B(_1385_),
    .A(net300),
    .Y(_1444_));
 sky130_as_sc_hs__buff_2 _3539_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1444_),
    .Y(_0105_));
 sky130_as_sc_hs__mux2_2 _3540_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1443_),
    .B(_1390_),
    .A(net356),
    .Y(_1445_));
 sky130_as_sc_hs__buff_2 _3541_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1445_),
    .Y(_0106_));
 sky130_as_sc_hs__mux2_2 _3542_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1443_),
    .B(_1392_),
    .A(net514),
    .Y(_1446_));
 sky130_as_sc_hs__buff_2 _3543_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1446_),
    .Y(_0107_));
 sky130_as_sc_hs__mux2_2 _3544_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1443_),
    .B(_1394_),
    .A(net411),
    .Y(_1447_));
 sky130_as_sc_hs__buff_2 _3545_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1447_),
    .Y(_0108_));
 sky130_as_sc_hs__mux2_2 _3546_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1443_),
    .B(_1396_),
    .A(net439),
    .Y(_1448_));
 sky130_as_sc_hs__buff_2 _3547_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1448_),
    .Y(_0109_));
 sky130_as_sc_hs__mux2_2 _3548_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1443_),
    .B(_1398_),
    .A(net414),
    .Y(_1449_));
 sky130_as_sc_hs__buff_2 _3549_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1449_),
    .Y(_0110_));
 sky130_as_sc_hs__buff_2 _3550_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1218_),
    .Y(_1450_));
 sky130_as_sc_hs__nor2_4 _3551_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1266_),
    .B(_1411_),
    .Y(_1451_));
 sky130_as_sc_hs__mux2_2 _3552_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1451_),
    .B(_1450_),
    .A(net497),
    .Y(_1452_));
 sky130_as_sc_hs__buff_2 _3553_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1452_),
    .Y(_0111_));
 sky130_as_sc_hs__buff_2 _3554_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1230_),
    .Y(_1453_));
 sky130_as_sc_hs__mux2_2 _3555_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1451_),
    .B(_1453_),
    .A(net510),
    .Y(_1454_));
 sky130_as_sc_hs__buff_2 _3556_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1454_),
    .Y(_0112_));
 sky130_as_sc_hs__buff_2 _3557_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1235_),
    .Y(_1455_));
 sky130_as_sc_hs__mux2_2 _3558_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1451_),
    .B(_1455_),
    .A(net336),
    .Y(_1456_));
 sky130_as_sc_hs__buff_2 _3559_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1456_),
    .Y(_0113_));
 sky130_as_sc_hs__buff_2 _3560_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1240_),
    .Y(_1457_));
 sky130_as_sc_hs__mux2_2 _3561_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1451_),
    .B(_1457_),
    .A(net541),
    .Y(_1458_));
 sky130_as_sc_hs__buff_2 _3562_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1458_),
    .Y(_0114_));
 sky130_as_sc_hs__buff_2 _3563_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1247_),
    .Y(_1459_));
 sky130_as_sc_hs__mux2_2 _3564_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1451_),
    .B(_1459_),
    .A(net507),
    .Y(_1460_));
 sky130_as_sc_hs__buff_2 _3565_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1460_),
    .Y(_0115_));
 sky130_as_sc_hs__buff_2 _3566_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1252_),
    .Y(_1461_));
 sky130_as_sc_hs__mux2_2 _3567_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1451_),
    .B(_1461_),
    .A(net242),
    .Y(_1462_));
 sky130_as_sc_hs__buff_2 _3568_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1462_),
    .Y(_0116_));
 sky130_as_sc_hs__nor2_4 _3569_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1256_),
    .B(_1276_),
    .Y(_1463_));
 sky130_as_sc_hs__mux2_2 _3570_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1463_),
    .B(_1450_),
    .A(net307),
    .Y(_1464_));
 sky130_as_sc_hs__buff_2 _3571_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1464_),
    .Y(_0117_));
 sky130_as_sc_hs__mux2_2 _3572_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1463_),
    .B(_1453_),
    .A(net357),
    .Y(_1465_));
 sky130_as_sc_hs__buff_2 _3573_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1465_),
    .Y(_0118_));
 sky130_as_sc_hs__mux2_2 _3574_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1463_),
    .B(_1455_),
    .A(net517),
    .Y(_1466_));
 sky130_as_sc_hs__buff_2 _3575_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1466_),
    .Y(_0119_));
 sky130_as_sc_hs__mux2_2 _3576_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1463_),
    .B(_1457_),
    .A(net329),
    .Y(_1467_));
 sky130_as_sc_hs__buff_2 _3577_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1467_),
    .Y(_0120_));
 sky130_as_sc_hs__mux2_2 _3578_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1463_),
    .B(_1459_),
    .A(net537),
    .Y(_1468_));
 sky130_as_sc_hs__buff_2 _3579_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1468_),
    .Y(_0121_));
 sky130_as_sc_hs__mux2_2 _3580_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1463_),
    .B(_1461_),
    .A(net546),
    .Y(_1469_));
 sky130_as_sc_hs__buff_2 _3581_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1469_),
    .Y(_0122_));
 sky130_as_sc_hs__clkbuff_4 _3582_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1217_),
    .Y(_1470_));
 sky130_as_sc_hs__or2_2 _3583_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0625_),
    .B(_1264_),
    .Y(_1471_));
 sky130_as_sc_hs__nor2_4 _3584_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1419_),
    .B(_1471_),
    .Y(_1472_));
 sky130_as_sc_hs__mux2_2 _3585_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1472_),
    .B(_1470_),
    .A(\RAM[58][0] ),
    .Y(_1473_));
 sky130_as_sc_hs__and2_2 _3586_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net146),
    .B(_1473_),
    .Y(_1474_));
 sky130_as_sc_hs__buff_2 _3587_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1474_),
    .Y(_0123_));
 sky130_as_sc_hs__buff_4 _3588_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1229_),
    .Y(_1475_));
 sky130_as_sc_hs__mux2_2 _3589_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1472_),
    .B(_1475_),
    .A(\RAM[58][1] ),
    .Y(_1476_));
 sky130_as_sc_hs__and2_2 _3590_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net146),
    .B(_1476_),
    .Y(_1477_));
 sky130_as_sc_hs__buff_2 _3591_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1477_),
    .Y(_0124_));
 sky130_as_sc_hs__buff_4 _3592_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1234_),
    .Y(_1478_));
 sky130_as_sc_hs__mux2_2 _3593_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1472_),
    .B(_1478_),
    .A(\RAM[58][2] ),
    .Y(_1479_));
 sky130_as_sc_hs__and2_2 _3594_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net146),
    .B(_1479_),
    .Y(_1480_));
 sky130_as_sc_hs__buff_2 _3595_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1480_),
    .Y(_0125_));
 sky130_as_sc_hs__buff_4 _3596_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1239_),
    .Y(_1481_));
 sky130_as_sc_hs__mux2_2 _3597_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1472_),
    .B(_1481_),
    .A(\RAM[58][3] ),
    .Y(_1482_));
 sky130_as_sc_hs__and2_2 _3598_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net146),
    .B(_1482_),
    .Y(_1483_));
 sky130_as_sc_hs__buff_2 _3599_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1483_),
    .Y(_0126_));
 sky130_as_sc_hs__buff_4 _3600_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1246_),
    .Y(_1484_));
 sky130_as_sc_hs__mux2_2 _3601_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1472_),
    .B(_1484_),
    .A(\RAM[58][4] ),
    .Y(_1485_));
 sky130_as_sc_hs__and2_2 _3602_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net146),
    .B(_1485_),
    .Y(_1486_));
 sky130_as_sc_hs__buff_2 _3603_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1486_),
    .Y(_0127_));
 sky130_as_sc_hs__buff_4 _3604_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1251_),
    .Y(_1487_));
 sky130_as_sc_hs__mux2_2 _3605_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1472_),
    .B(_1487_),
    .A(\RAM[58][5] ),
    .Y(_1488_));
 sky130_as_sc_hs__and2_2 _3606_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net146),
    .B(_1488_),
    .Y(_1489_));
 sky130_as_sc_hs__buff_2 _3607_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1489_),
    .Y(_0128_));
 sky130_as_sc_hs__clkbuff_11 _3608_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1471_),
    .Y(_1490_));
 sky130_as_sc_hs__nor2_4 _3609_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1225_),
    .B(_1490_),
    .Y(_1491_));
 sky130_as_sc_hs__mux2_2 _3610_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1491_),
    .B(_1450_),
    .A(net475),
    .Y(_1492_));
 sky130_as_sc_hs__buff_2 _3611_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1492_),
    .Y(_0129_));
 sky130_as_sc_hs__mux2_2 _3612_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1491_),
    .B(_1453_),
    .A(net524),
    .Y(_1493_));
 sky130_as_sc_hs__buff_2 _3613_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1493_),
    .Y(_0130_));
 sky130_as_sc_hs__mux2_2 _3614_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1491_),
    .B(_1455_),
    .A(net538),
    .Y(_1494_));
 sky130_as_sc_hs__buff_2 _3615_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1494_),
    .Y(_0131_));
 sky130_as_sc_hs__mux2_2 _3616_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1491_),
    .B(_1457_),
    .A(net479),
    .Y(_1495_));
 sky130_as_sc_hs__buff_2 _3617_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1495_),
    .Y(_0132_));
 sky130_as_sc_hs__mux2_2 _3618_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1491_),
    .B(_1459_),
    .A(net298),
    .Y(_1496_));
 sky130_as_sc_hs__buff_2 _3619_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1496_),
    .Y(_0133_));
 sky130_as_sc_hs__mux2_2 _3620_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1491_),
    .B(_1461_),
    .A(net235),
    .Y(_1497_));
 sky130_as_sc_hs__buff_2 _3621_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1497_),
    .Y(_0134_));
 sky130_as_sc_hs__nor2_4 _3622_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1225_),
    .B(_1402_),
    .Y(_1498_));
 sky130_as_sc_hs__mux2_2 _3623_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1498_),
    .B(_1450_),
    .A(net255),
    .Y(_1499_));
 sky130_as_sc_hs__buff_2 _3624_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1499_),
    .Y(_0135_));
 sky130_as_sc_hs__mux2_2 _3625_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1498_),
    .B(_1453_),
    .A(net316),
    .Y(_1500_));
 sky130_as_sc_hs__buff_2 _3626_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1500_),
    .Y(_0136_));
 sky130_as_sc_hs__mux2_2 _3627_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1498_),
    .B(_1455_),
    .A(net335),
    .Y(_1501_));
 sky130_as_sc_hs__buff_2 _3628_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1501_),
    .Y(_0137_));
 sky130_as_sc_hs__mux2_2 _3629_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1498_),
    .B(_1457_),
    .A(net281),
    .Y(_1502_));
 sky130_as_sc_hs__buff_2 _3630_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1502_),
    .Y(_0138_));
 sky130_as_sc_hs__mux2_2 _3631_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1498_),
    .B(_1459_),
    .A(net243),
    .Y(_1503_));
 sky130_as_sc_hs__buff_2 _3632_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1503_),
    .Y(_0139_));
 sky130_as_sc_hs__mux2_2 _3633_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1498_),
    .B(_1461_),
    .A(net312),
    .Y(_1504_));
 sky130_as_sc_hs__buff_2 _3634_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1504_),
    .Y(_0140_));
 sky130_as_sc_hs__nor2_4 _3635_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1223_),
    .B(_1276_),
    .Y(_1505_));
 sky130_as_sc_hs__mux2_2 _3636_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1505_),
    .B(_1450_),
    .A(net295),
    .Y(_1506_));
 sky130_as_sc_hs__buff_2 _3637_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1506_),
    .Y(_0141_));
 sky130_as_sc_hs__mux2_2 _3638_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1505_),
    .B(_1453_),
    .A(net380),
    .Y(_1507_));
 sky130_as_sc_hs__buff_2 _3639_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1507_),
    .Y(_0142_));
 sky130_as_sc_hs__mux2_2 _3640_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1505_),
    .B(_1455_),
    .A(net350),
    .Y(_1508_));
 sky130_as_sc_hs__buff_2 _3641_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1508_),
    .Y(_0143_));
 sky130_as_sc_hs__mux2_2 _3642_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1505_),
    .B(_1457_),
    .A(net474),
    .Y(_1509_));
 sky130_as_sc_hs__buff_2 _3643_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1509_),
    .Y(_0144_));
 sky130_as_sc_hs__mux2_2 _3644_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1505_),
    .B(_1459_),
    .A(net327),
    .Y(_1510_));
 sky130_as_sc_hs__buff_2 _3645_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1510_),
    .Y(_0145_));
 sky130_as_sc_hs__mux2_2 _3646_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1505_),
    .B(_1461_),
    .A(net545),
    .Y(_1511_));
 sky130_as_sc_hs__buff_2 _3647_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1511_),
    .Y(_0146_));
 sky130_as_sc_hs__nor2_4 _3648_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1400_),
    .B(_1366_),
    .Y(_1512_));
 sky130_as_sc_hs__mux2_2 _3649_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1512_),
    .B(_1450_),
    .A(net376),
    .Y(_1513_));
 sky130_as_sc_hs__buff_2 _3650_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1513_),
    .Y(_0147_));
 sky130_as_sc_hs__mux2_2 _3651_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1512_),
    .B(_1453_),
    .A(net488),
    .Y(_1514_));
 sky130_as_sc_hs__buff_2 _3652_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1514_),
    .Y(_0148_));
 sky130_as_sc_hs__mux2_2 _3653_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1512_),
    .B(_1455_),
    .A(net388),
    .Y(_1515_));
 sky130_as_sc_hs__buff_2 _3654_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1515_),
    .Y(_0149_));
 sky130_as_sc_hs__mux2_2 _3655_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1512_),
    .B(_1457_),
    .A(net261),
    .Y(_1516_));
 sky130_as_sc_hs__buff_2 _3656_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1516_),
    .Y(_0150_));
 sky130_as_sc_hs__mux2_2 _3657_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1512_),
    .B(_1459_),
    .A(net489),
    .Y(_1517_));
 sky130_as_sc_hs__buff_2 _3658_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1517_),
    .Y(_0151_));
 sky130_as_sc_hs__mux2_2 _3659_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1512_),
    .B(_1461_),
    .A(net365),
    .Y(_1518_));
 sky130_as_sc_hs__buff_2 _3660_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1518_),
    .Y(_0152_));
 sky130_as_sc_hs__nor2_4 _3661_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1225_),
    .B(_1275_),
    .Y(_1519_));
 sky130_as_sc_hs__mux2_2 _3662_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1519_),
    .B(_1450_),
    .A(net554),
    .Y(_1520_));
 sky130_as_sc_hs__buff_2 _3663_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1520_),
    .Y(_0153_));
 sky130_as_sc_hs__mux2_2 _3664_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1519_),
    .B(_1453_),
    .A(net522),
    .Y(_1521_));
 sky130_as_sc_hs__buff_2 _3665_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1521_),
    .Y(_0154_));
 sky130_as_sc_hs__mux2_2 _3666_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1519_),
    .B(_1455_),
    .A(net567),
    .Y(_1522_));
 sky130_as_sc_hs__buff_2 _3667_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1522_),
    .Y(_0155_));
 sky130_as_sc_hs__mux2_2 _3668_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1519_),
    .B(_1457_),
    .A(net484),
    .Y(_1523_));
 sky130_as_sc_hs__buff_2 _3669_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1523_),
    .Y(_0156_));
 sky130_as_sc_hs__mux2_2 _3670_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1519_),
    .B(_1459_),
    .A(net314),
    .Y(_1524_));
 sky130_as_sc_hs__buff_2 _3671_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1524_),
    .Y(_0157_));
 sky130_as_sc_hs__mux2_2 _3672_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1519_),
    .B(_1461_),
    .A(net288),
    .Y(_1525_));
 sky130_as_sc_hs__buff_2 _3673_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1525_),
    .Y(_0158_));
 sky130_as_sc_hs__clkbuff_4 _3674_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1218_),
    .Y(_1526_));
 sky130_as_sc_hs__nor2_4 _3675_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1366_),
    .B(_1428_),
    .Y(_1527_));
 sky130_as_sc_hs__mux2_2 _3676_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1527_),
    .B(_1526_),
    .A(net551),
    .Y(_1528_));
 sky130_as_sc_hs__buff_2 _3677_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1528_),
    .Y(_0159_));
 sky130_as_sc_hs__clkbuff_4 _3678_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1230_),
    .Y(_1529_));
 sky130_as_sc_hs__mux2_2 _3679_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1527_),
    .B(_1529_),
    .A(net562),
    .Y(_1530_));
 sky130_as_sc_hs__buff_2 _3680_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1530_),
    .Y(_0160_));
 sky130_as_sc_hs__clkbuff_4 _3681_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1235_),
    .Y(_1531_));
 sky130_as_sc_hs__mux2_2 _3682_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1527_),
    .B(_1531_),
    .A(net233),
    .Y(_1532_));
 sky130_as_sc_hs__buff_2 _3683_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1532_),
    .Y(_0161_));
 sky130_as_sc_hs__clkbuff_4 _3684_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1240_),
    .Y(_1533_));
 sky130_as_sc_hs__mux2_2 _3685_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1527_),
    .B(_1533_),
    .A(net472),
    .Y(_1534_));
 sky130_as_sc_hs__buff_2 _3686_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1534_),
    .Y(_0162_));
 sky130_as_sc_hs__buff_4 _3687_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1247_),
    .Y(_1535_));
 sky130_as_sc_hs__mux2_2 _3688_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1527_),
    .B(_1535_),
    .A(net278),
    .Y(_1536_));
 sky130_as_sc_hs__buff_2 _3689_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1536_),
    .Y(_0163_));
 sky130_as_sc_hs__buff_4 _3690_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1252_),
    .Y(_1537_));
 sky130_as_sc_hs__mux2_2 _3691_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1527_),
    .B(_1537_),
    .A(net237),
    .Y(_1538_));
 sky130_as_sc_hs__buff_2 _3692_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1538_),
    .Y(_0164_));
 sky130_as_sc_hs__nor2_4 _3693_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1256_),
    .B(_1369_),
    .Y(_1539_));
 sky130_as_sc_hs__mux2_2 _3694_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1539_),
    .B(_1526_),
    .A(net337),
    .Y(_1540_));
 sky130_as_sc_hs__buff_2 _3695_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1540_),
    .Y(_0165_));
 sky130_as_sc_hs__mux2_2 _3696_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1539_),
    .B(_1529_),
    .A(net378),
    .Y(_1541_));
 sky130_as_sc_hs__buff_2 _3697_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1541_),
    .Y(_0166_));
 sky130_as_sc_hs__mux2_2 _3698_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1539_),
    .B(_1531_),
    .A(net490),
    .Y(_1542_));
 sky130_as_sc_hs__buff_2 _3699_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1542_),
    .Y(_0167_));
 sky130_as_sc_hs__mux2_2 _3700_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1539_),
    .B(_1533_),
    .A(net239),
    .Y(_1543_));
 sky130_as_sc_hs__buff_2 _3701_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1543_),
    .Y(_0168_));
 sky130_as_sc_hs__mux2_2 _3702_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1539_),
    .B(_1535_),
    .A(net308),
    .Y(_1544_));
 sky130_as_sc_hs__buff_2 _3703_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1544_),
    .Y(_0169_));
 sky130_as_sc_hs__mux2_2 _3704_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1539_),
    .B(_1537_),
    .A(net383),
    .Y(_1545_));
 sky130_as_sc_hs__buff_2 _3705_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1545_),
    .Y(_0170_));
 sky130_as_sc_hs__nor2_4 _3706_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1400_),
    .B(_1490_),
    .Y(_1546_));
 sky130_as_sc_hs__mux2_2 _3707_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1546_),
    .B(_1526_),
    .A(net420),
    .Y(_1547_));
 sky130_as_sc_hs__buff_2 _3708_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1547_),
    .Y(_0171_));
 sky130_as_sc_hs__mux2_2 _3709_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1546_),
    .B(_1529_),
    .A(net450),
    .Y(_1548_));
 sky130_as_sc_hs__buff_2 _3710_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1548_),
    .Y(_0172_));
 sky130_as_sc_hs__mux2_2 _3711_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1546_),
    .B(_1531_),
    .A(net508),
    .Y(_1549_));
 sky130_as_sc_hs__buff_2 _3712_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1549_),
    .Y(_0173_));
 sky130_as_sc_hs__mux2_2 _3713_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1546_),
    .B(_1533_),
    .A(net539),
    .Y(_1550_));
 sky130_as_sc_hs__buff_2 _3714_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1550_),
    .Y(_0174_));
 sky130_as_sc_hs__mux2_2 _3715_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1546_),
    .B(_1535_),
    .A(net552),
    .Y(_1551_));
 sky130_as_sc_hs__buff_2 _3716_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1551_),
    .Y(_0175_));
 sky130_as_sc_hs__mux2_2 _3717_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1546_),
    .B(_1537_),
    .A(net495),
    .Y(_1552_));
 sky130_as_sc_hs__buff_2 _3718_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1552_),
    .Y(_0176_));
 sky130_as_sc_hs__or2_2 _3719_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0631_),
    .B(_1367_),
    .Y(_1553_));
 sky130_as_sc_hs__buff_6 _3720_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1553_),
    .Y(_1554_));
 sky130_as_sc_hs__nor2_4 _3721_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1266_),
    .B(_1554_),
    .Y(_1555_));
 sky130_as_sc_hs__mux2_2 _3722_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1555_),
    .B(_1526_),
    .A(net254),
    .Y(_1556_));
 sky130_as_sc_hs__buff_2 _3723_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1556_),
    .Y(_0177_));
 sky130_as_sc_hs__mux2_2 _3724_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1555_),
    .B(_1529_),
    .A(net387),
    .Y(_1557_));
 sky130_as_sc_hs__buff_2 _3725_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1557_),
    .Y(_0178_));
 sky130_as_sc_hs__mux2_2 _3726_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1555_),
    .B(_1531_),
    .A(net499),
    .Y(_1558_));
 sky130_as_sc_hs__buff_2 _3727_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1558_),
    .Y(_0179_));
 sky130_as_sc_hs__mux2_2 _3728_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1555_),
    .B(_1533_),
    .A(net210),
    .Y(_1559_));
 sky130_as_sc_hs__buff_2 _3729_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1559_),
    .Y(_0180_));
 sky130_as_sc_hs__mux2_2 _3730_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1555_),
    .B(_1535_),
    .A(net432),
    .Y(_1560_));
 sky130_as_sc_hs__buff_2 _3731_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1560_),
    .Y(_0181_));
 sky130_as_sc_hs__mux2_2 _3732_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1555_),
    .B(_1537_),
    .A(net360),
    .Y(_1561_));
 sky130_as_sc_hs__buff_2 _3733_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1561_),
    .Y(_0182_));
 sky130_as_sc_hs__nor2_4 _3734_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1256_),
    .B(_1411_),
    .Y(_1562_));
 sky130_as_sc_hs__mux2_2 _3735_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1562_),
    .B(_1526_),
    .A(net323),
    .Y(_1563_));
 sky130_as_sc_hs__buff_2 _3736_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1563_),
    .Y(_0183_));
 sky130_as_sc_hs__mux2_2 _3737_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1562_),
    .B(_1529_),
    .A(net302),
    .Y(_1564_));
 sky130_as_sc_hs__buff_2 _3738_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1564_),
    .Y(_0184_));
 sky130_as_sc_hs__mux2_2 _3739_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1562_),
    .B(_1531_),
    .A(net309),
    .Y(_1565_));
 sky130_as_sc_hs__buff_2 _3740_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1565_),
    .Y(_0185_));
 sky130_as_sc_hs__mux2_2 _3741_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1562_),
    .B(_1533_),
    .A(net466),
    .Y(_1566_));
 sky130_as_sc_hs__buff_2 _3742_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1566_),
    .Y(_0186_));
 sky130_as_sc_hs__mux2_2 _3743_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1562_),
    .B(_1535_),
    .A(net321),
    .Y(_1567_));
 sky130_as_sc_hs__buff_2 _3744_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1567_),
    .Y(_0187_));
 sky130_as_sc_hs__mux2_2 _3745_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1562_),
    .B(_1537_),
    .A(net285),
    .Y(_1568_));
 sky130_as_sc_hs__buff_2 _3746_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1568_),
    .Y(_0188_));
 sky130_as_sc_hs__aoi31_2 _3747_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net101),
    .B(_0695_),
    .C(_1213_),
    .D(_1156_),
    .Y(_1569_));
 sky130_as_sc_hs__nor2_4 _3748_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1553_),
    .B(_1569_),
    .Y(_1570_));
 sky130_as_sc_hs__mux2_2 _3749_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1570_),
    .B(_1526_),
    .A(net305),
    .Y(_1571_));
 sky130_as_sc_hs__buff_2 _3750_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1571_),
    .Y(_0189_));
 sky130_as_sc_hs__mux2_2 _3751_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1570_),
    .B(_1529_),
    .A(net529),
    .Y(_1572_));
 sky130_as_sc_hs__buff_2 _3752_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1572_),
    .Y(_0190_));
 sky130_as_sc_hs__mux2_2 _3753_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1570_),
    .B(_1531_),
    .A(net266),
    .Y(_1573_));
 sky130_as_sc_hs__buff_2 _3754_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1573_),
    .Y(_0191_));
 sky130_as_sc_hs__mux2_2 _3755_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1570_),
    .B(_1533_),
    .A(net274),
    .Y(_1574_));
 sky130_as_sc_hs__buff_2 _3756_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1574_),
    .Y(_0192_));
 sky130_as_sc_hs__mux2_2 _3757_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1570_),
    .B(_1535_),
    .A(net292),
    .Y(_1575_));
 sky130_as_sc_hs__buff_2 _3758_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1575_),
    .Y(_0193_));
 sky130_as_sc_hs__mux2_2 _3759_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1570_),
    .B(_1537_),
    .A(net359),
    .Y(_1576_));
 sky130_as_sc_hs__buff_2 _3760_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1576_),
    .Y(_0194_));
 sky130_as_sc_hs__nor2_4 _3761_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1223_),
    .B(_1411_),
    .Y(_1577_));
 sky130_as_sc_hs__mux2_2 _3762_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1577_),
    .B(_1526_),
    .A(net225),
    .Y(_1578_));
 sky130_as_sc_hs__buff_2 _3763_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1578_),
    .Y(_0195_));
 sky130_as_sc_hs__mux2_2 _3764_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1577_),
    .B(_1529_),
    .A(net303),
    .Y(_1579_));
 sky130_as_sc_hs__buff_2 _3765_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1579_),
    .Y(_0196_));
 sky130_as_sc_hs__mux2_2 _3766_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1577_),
    .B(_1531_),
    .A(net381),
    .Y(_1580_));
 sky130_as_sc_hs__buff_2 _3767_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1580_),
    .Y(_0197_));
 sky130_as_sc_hs__mux2_2 _3768_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1577_),
    .B(_1533_),
    .A(net548),
    .Y(_1581_));
 sky130_as_sc_hs__buff_2 _3769_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1581_),
    .Y(_0198_));
 sky130_as_sc_hs__mux2_2 _3770_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1577_),
    .B(_1535_),
    .A(net428),
    .Y(_1582_));
 sky130_as_sc_hs__buff_2 _3771_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1582_),
    .Y(_0199_));
 sky130_as_sc_hs__mux2_2 _3772_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1577_),
    .B(_1537_),
    .A(net223),
    .Y(_1583_));
 sky130_as_sc_hs__buff_2 _3773_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1583_),
    .Y(_0200_));
 sky130_as_sc_hs__clkbuff_4 _3774_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1218_),
    .Y(_1584_));
 sky130_as_sc_hs__nor2_4 _3775_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1369_),
    .B(_1402_),
    .Y(_1585_));
 sky130_as_sc_hs__mux2_2 _3776_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1585_),
    .B(_1584_),
    .A(net196),
    .Y(_1586_));
 sky130_as_sc_hs__buff_2 _3777_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1586_),
    .Y(_0201_));
 sky130_as_sc_hs__buff_2 _3778_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1230_),
    .Y(_1587_));
 sky130_as_sc_hs__mux2_2 _3779_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1585_),
    .B(_1587_),
    .A(net273),
    .Y(_1588_));
 sky130_as_sc_hs__buff_2 _3780_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1588_),
    .Y(_0202_));
 sky130_as_sc_hs__buff_2 _3781_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1235_),
    .Y(_1589_));
 sky130_as_sc_hs__mux2_2 _3782_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1585_),
    .B(_1589_),
    .A(net453),
    .Y(_1590_));
 sky130_as_sc_hs__buff_2 _3783_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1590_),
    .Y(_0203_));
 sky130_as_sc_hs__buff_2 _3784_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1240_),
    .Y(_1591_));
 sky130_as_sc_hs__mux2_2 _3785_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1585_),
    .B(_1591_),
    .A(net465),
    .Y(_1592_));
 sky130_as_sc_hs__buff_2 _3786_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1592_),
    .Y(_0204_));
 sky130_as_sc_hs__buff_2 _3787_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1247_),
    .Y(_1593_));
 sky130_as_sc_hs__mux2_2 _3788_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1585_),
    .B(_1593_),
    .A(net559),
    .Y(_1594_));
 sky130_as_sc_hs__buff_2 _3789_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1594_),
    .Y(_0205_));
 sky130_as_sc_hs__buff_2 _3790_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1252_),
    .Y(_1595_));
 sky130_as_sc_hs__mux2_2 _3791_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1585_),
    .B(_1595_),
    .A(net444),
    .Y(_1596_));
 sky130_as_sc_hs__buff_2 _3792_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1596_),
    .Y(_0206_));
 sky130_as_sc_hs__nor2_4 _3793_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1366_),
    .B(_1411_),
    .Y(_1597_));
 sky130_as_sc_hs__mux2_2 _3794_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1597_),
    .B(_1584_),
    .A(net291),
    .Y(_1598_));
 sky130_as_sc_hs__buff_2 _3795_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1598_),
    .Y(_0207_));
 sky130_as_sc_hs__mux2_2 _3796_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1597_),
    .B(_1587_),
    .A(net260),
    .Y(_1599_));
 sky130_as_sc_hs__buff_2 _3797_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1599_),
    .Y(_0208_));
 sky130_as_sc_hs__mux2_2 _3798_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1597_),
    .B(_1589_),
    .A(net313),
    .Y(_1600_));
 sky130_as_sc_hs__buff_2 _3799_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1600_),
    .Y(_0209_));
 sky130_as_sc_hs__mux2_2 _3800_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1597_),
    .B(_1591_),
    .A(net389),
    .Y(_1601_));
 sky130_as_sc_hs__buff_2 _3801_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1601_),
    .Y(_0210_));
 sky130_as_sc_hs__mux2_2 _3802_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1597_),
    .B(_1593_),
    .A(net361),
    .Y(_1602_));
 sky130_as_sc_hs__buff_2 _3803_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1602_),
    .Y(_0211_));
 sky130_as_sc_hs__mux2_2 _3804_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1597_),
    .B(_1595_),
    .A(net476),
    .Y(_1603_));
 sky130_as_sc_hs__buff_2 _3805_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1603_),
    .Y(_0212_));
 sky130_as_sc_hs__nor2_4 _3806_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1275_),
    .B(_1369_),
    .Y(_1604_));
 sky130_as_sc_hs__mux2_2 _3807_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1604_),
    .B(_1584_),
    .A(net318),
    .Y(_1605_));
 sky130_as_sc_hs__buff_2 _3808_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1605_),
    .Y(_0213_));
 sky130_as_sc_hs__mux2_2 _3809_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1604_),
    .B(_1587_),
    .A(net399),
    .Y(_1606_));
 sky130_as_sc_hs__buff_2 _3810_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1606_),
    .Y(_0214_));
 sky130_as_sc_hs__mux2_2 _3811_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1604_),
    .B(_1589_),
    .A(net297),
    .Y(_1607_));
 sky130_as_sc_hs__buff_2 _3812_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1607_),
    .Y(_0215_));
 sky130_as_sc_hs__mux2_2 _3813_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1604_),
    .B(_1591_),
    .A(net330),
    .Y(_1608_));
 sky130_as_sc_hs__buff_2 _3814_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1608_),
    .Y(_0216_));
 sky130_as_sc_hs__mux2_2 _3815_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1604_),
    .B(_1593_),
    .A(net568),
    .Y(_1609_));
 sky130_as_sc_hs__buff_2 _3816_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1609_),
    .Y(_0217_));
 sky130_as_sc_hs__mux2_2 _3817_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1604_),
    .B(_1595_),
    .A(net478),
    .Y(_1610_));
 sky130_as_sc_hs__buff_2 _3818_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1610_),
    .Y(_0218_));
 sky130_as_sc_hs__nor2_4 _3819_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1410_),
    .B(_1490_),
    .Y(_1611_));
 sky130_as_sc_hs__mux2_2 _3820_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1611_),
    .B(_1584_),
    .A(net207),
    .Y(_1612_));
 sky130_as_sc_hs__buff_2 _3821_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1612_),
    .Y(_0219_));
 sky130_as_sc_hs__mux2_2 _3822_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1611_),
    .B(_1587_),
    .A(net390),
    .Y(_1613_));
 sky130_as_sc_hs__buff_2 _3823_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1613_),
    .Y(_0220_));
 sky130_as_sc_hs__mux2_2 _3824_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1611_),
    .B(_1589_),
    .A(net442),
    .Y(_1614_));
 sky130_as_sc_hs__buff_2 _3825_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1614_),
    .Y(_0221_));
 sky130_as_sc_hs__mux2_2 _3826_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1611_),
    .B(_1591_),
    .A(net248),
    .Y(_1615_));
 sky130_as_sc_hs__buff_2 _3827_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1615_),
    .Y(_0222_));
 sky130_as_sc_hs__mux2_2 _3828_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1611_),
    .B(_1593_),
    .A(net496),
    .Y(_1616_));
 sky130_as_sc_hs__buff_2 _3829_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1616_),
    .Y(_0223_));
 sky130_as_sc_hs__mux2_2 _3830_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1611_),
    .B(_1595_),
    .A(net511),
    .Y(_1617_));
 sky130_as_sc_hs__buff_2 _3831_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1617_),
    .Y(_0224_));
 sky130_as_sc_hs__nor2_4 _3832_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1369_),
    .B(_1490_),
    .Y(_1618_));
 sky130_as_sc_hs__mux2_2 _3833_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1618_),
    .B(_1584_),
    .A(net211),
    .Y(_1619_));
 sky130_as_sc_hs__buff_2 _3834_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1619_),
    .Y(_0225_));
 sky130_as_sc_hs__mux2_2 _3835_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1618_),
    .B(_1587_),
    .A(net251),
    .Y(_1620_));
 sky130_as_sc_hs__buff_2 _3836_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1620_),
    .Y(_0226_));
 sky130_as_sc_hs__mux2_2 _3837_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1618_),
    .B(_1589_),
    .A(net504),
    .Y(_1621_));
 sky130_as_sc_hs__buff_2 _3838_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1621_),
    .Y(_0227_));
 sky130_as_sc_hs__mux2_2 _3839_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1618_),
    .B(_1591_),
    .A(net519),
    .Y(_1622_));
 sky130_as_sc_hs__buff_2 _3840_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1622_),
    .Y(_0228_));
 sky130_as_sc_hs__mux2_2 _3841_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1618_),
    .B(_1593_),
    .A(net557),
    .Y(_1623_));
 sky130_as_sc_hs__buff_2 _3842_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1623_),
    .Y(_0229_));
 sky130_as_sc_hs__mux2_2 _3843_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1618_),
    .B(_1595_),
    .A(net382),
    .Y(_1624_));
 sky130_as_sc_hs__buff_2 _3844_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1624_),
    .Y(_0230_));
 sky130_as_sc_hs__nor2_4 _3845_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1275_),
    .B(_1411_),
    .Y(_1625_));
 sky130_as_sc_hs__mux2_2 _3846_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1625_),
    .B(_1584_),
    .A(net319),
    .Y(_1626_));
 sky130_as_sc_hs__buff_2 _3847_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1626_),
    .Y(_0231_));
 sky130_as_sc_hs__mux2_2 _3848_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1625_),
    .B(_1587_),
    .A(net226),
    .Y(_1627_));
 sky130_as_sc_hs__buff_2 _3849_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1627_),
    .Y(_0232_));
 sky130_as_sc_hs__mux2_2 _3850_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1625_),
    .B(_1589_),
    .A(net247),
    .Y(_1628_));
 sky130_as_sc_hs__buff_2 _3851_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1628_),
    .Y(_0233_));
 sky130_as_sc_hs__mux2_2 _3852_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1625_),
    .B(_1591_),
    .A(net447),
    .Y(_1629_));
 sky130_as_sc_hs__buff_2 _3853_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1629_),
    .Y(_0234_));
 sky130_as_sc_hs__mux2_2 _3854_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1625_),
    .B(_1593_),
    .A(net289),
    .Y(_1630_));
 sky130_as_sc_hs__buff_2 _3855_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1630_),
    .Y(_0235_));
 sky130_as_sc_hs__mux2_2 _3856_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1625_),
    .B(_1595_),
    .A(net262),
    .Y(_1631_));
 sky130_as_sc_hs__buff_2 _3857_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1631_),
    .Y(_0236_));
 sky130_as_sc_hs__nor2_4 _3858_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1275_),
    .B(_1428_),
    .Y(_1632_));
 sky130_as_sc_hs__mux2_2 _3859_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1632_),
    .B(_1584_),
    .A(net470),
    .Y(_1633_));
 sky130_as_sc_hs__buff_2 _3860_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1633_),
    .Y(_0237_));
 sky130_as_sc_hs__mux2_2 _3861_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1632_),
    .B(_1587_),
    .A(net464),
    .Y(_1634_));
 sky130_as_sc_hs__buff_2 _3862_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1634_),
    .Y(_0238_));
 sky130_as_sc_hs__mux2_2 _3863_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1632_),
    .B(_1589_),
    .A(net563),
    .Y(_1635_));
 sky130_as_sc_hs__buff_2 _3864_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1635_),
    .Y(_0239_));
 sky130_as_sc_hs__mux2_2 _3865_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1632_),
    .B(_1591_),
    .A(net569),
    .Y(_1636_));
 sky130_as_sc_hs__buff_2 _3866_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1636_),
    .Y(_0240_));
 sky130_as_sc_hs__mux2_2 _3867_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1632_),
    .B(_1593_),
    .A(net341),
    .Y(_1637_));
 sky130_as_sc_hs__buff_2 _3868_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1637_),
    .Y(_0241_));
 sky130_as_sc_hs__mux2_2 _3869_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1632_),
    .B(_1595_),
    .A(net486),
    .Y(_1638_));
 sky130_as_sc_hs__buff_2 _3870_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1638_),
    .Y(_0242_));
 sky130_as_sc_hs__buff_4 _3871_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1218_),
    .Y(_1639_));
 sky130_as_sc_hs__nor2_4 _3872_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1402_),
    .B(_1411_),
    .Y(_1640_));
 sky130_as_sc_hs__mux2_2 _3873_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1640_),
    .B(_1639_),
    .A(net373),
    .Y(_1641_));
 sky130_as_sc_hs__buff_2 _3874_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1641_),
    .Y(_0243_));
 sky130_as_sc_hs__buff_4 _3875_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1230_),
    .Y(_1642_));
 sky130_as_sc_hs__mux2_2 _3876_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1640_),
    .B(_1642_),
    .A(net485),
    .Y(_1643_));
 sky130_as_sc_hs__buff_2 _3877_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1643_),
    .Y(_0244_));
 sky130_as_sc_hs__buff_4 _3878_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1235_),
    .Y(_1644_));
 sky130_as_sc_hs__mux2_2 _3879_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1640_),
    .B(_1644_),
    .A(net197),
    .Y(_1645_));
 sky130_as_sc_hs__buff_2 _3880_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1645_),
    .Y(_0245_));
 sky130_as_sc_hs__buff_4 _3881_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1240_),
    .Y(_1646_));
 sky130_as_sc_hs__mux2_2 _3882_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1640_),
    .B(_1646_),
    .A(net252),
    .Y(_1647_));
 sky130_as_sc_hs__buff_2 _3883_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1647_),
    .Y(_0246_));
 sky130_as_sc_hs__buff_4 _3884_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1247_),
    .Y(_1648_));
 sky130_as_sc_hs__mux2_2 _3885_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1640_),
    .B(_1648_),
    .A(net536),
    .Y(_1649_));
 sky130_as_sc_hs__buff_2 _3886_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1649_),
    .Y(_0247_));
 sky130_as_sc_hs__buff_4 _3887_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1252_),
    .Y(_1650_));
 sky130_as_sc_hs__mux2_2 _3888_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1640_),
    .B(_1650_),
    .A(net513),
    .Y(_1651_));
 sky130_as_sc_hs__buff_2 _3889_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1651_),
    .Y(_0248_));
 sky130_as_sc_hs__nor2_4 _3890_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1223_),
    .B(_1369_),
    .Y(_1652_));
 sky130_as_sc_hs__mux2_2 _3891_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1652_),
    .B(_1639_),
    .A(net208),
    .Y(_1653_));
 sky130_as_sc_hs__buff_2 _3892_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1653_),
    .Y(_0249_));
 sky130_as_sc_hs__mux2_2 _3893_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1652_),
    .B(_1642_),
    .A(net364),
    .Y(_1654_));
 sky130_as_sc_hs__buff_2 _3894_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1654_),
    .Y(_0250_));
 sky130_as_sc_hs__mux2_2 _3895_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1652_),
    .B(_1644_),
    .A(net440),
    .Y(_1655_));
 sky130_as_sc_hs__buff_2 _3896_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1655_),
    .Y(_0251_));
 sky130_as_sc_hs__mux2_2 _3897_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1652_),
    .B(_1646_),
    .A(net234),
    .Y(_1656_));
 sky130_as_sc_hs__buff_2 _3898_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1656_),
    .Y(_0252_));
 sky130_as_sc_hs__mux2_2 _3899_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1652_),
    .B(_1648_),
    .A(net340),
    .Y(_1657_));
 sky130_as_sc_hs__buff_2 _3900_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1657_),
    .Y(_0253_));
 sky130_as_sc_hs__mux2_2 _3901_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1652_),
    .B(_1650_),
    .A(net348),
    .Y(_1658_));
 sky130_as_sc_hs__buff_2 _3902_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1658_),
    .Y(_0254_));
 sky130_as_sc_hs__nor2_4 _3903_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1377_),
    .B(_1387_),
    .Y(_1659_));
 sky130_as_sc_hs__mux2_2 _3904_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1659_),
    .B(_1639_),
    .A(net232),
    .Y(_1660_));
 sky130_as_sc_hs__buff_2 _3905_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1660_),
    .Y(_0255_));
 sky130_as_sc_hs__mux2_2 _3906_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1659_),
    .B(_1642_),
    .A(net216),
    .Y(_1661_));
 sky130_as_sc_hs__buff_2 _3907_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1661_),
    .Y(_0256_));
 sky130_as_sc_hs__mux2_2 _3908_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1659_),
    .B(_1644_),
    .A(net438),
    .Y(_1662_));
 sky130_as_sc_hs__buff_2 _3909_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1662_),
    .Y(_0257_));
 sky130_as_sc_hs__mux2_2 _3910_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1659_),
    .B(_1646_),
    .A(net299),
    .Y(_1663_));
 sky130_as_sc_hs__buff_2 _3911_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1663_),
    .Y(_0258_));
 sky130_as_sc_hs__mux2_2 _3912_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1659_),
    .B(_1648_),
    .A(net306),
    .Y(_1664_));
 sky130_as_sc_hs__buff_2 _3913_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1664_),
    .Y(_0259_));
 sky130_as_sc_hs__mux2_2 _3914_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1659_),
    .B(_1650_),
    .A(net530),
    .Y(_1665_));
 sky130_as_sc_hs__buff_2 _3915_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1665_),
    .Y(_0260_));
 sky130_as_sc_hs__nor2_4 _3916_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1266_),
    .B(_1387_),
    .Y(_1666_));
 sky130_as_sc_hs__mux2_2 _3917_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1666_),
    .B(_1639_),
    .A(net230),
    .Y(_1667_));
 sky130_as_sc_hs__buff_2 _3918_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1667_),
    .Y(_0261_));
 sky130_as_sc_hs__mux2_2 _3919_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1666_),
    .B(_1642_),
    .A(net263),
    .Y(_1668_));
 sky130_as_sc_hs__buff_2 _3920_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1668_),
    .Y(_0262_));
 sky130_as_sc_hs__mux2_2 _3921_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1666_),
    .B(_1644_),
    .A(net218),
    .Y(_1669_));
 sky130_as_sc_hs__buff_2 _3922_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1669_),
    .Y(_0263_));
 sky130_as_sc_hs__mux2_2 _3923_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1666_),
    .B(_1646_),
    .A(net535),
    .Y(_1670_));
 sky130_as_sc_hs__buff_2 _3924_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1670_),
    .Y(_0264_));
 sky130_as_sc_hs__mux2_2 _3925_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1666_),
    .B(_1648_),
    .A(net282),
    .Y(_1671_));
 sky130_as_sc_hs__buff_2 _3926_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1671_),
    .Y(_0265_));
 sky130_as_sc_hs__mux2_2 _3927_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1666_),
    .B(_1650_),
    .A(net555),
    .Y(_1672_));
 sky130_as_sc_hs__buff_2 _3928_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1672_),
    .Y(_0266_));
 sky130_as_sc_hs__nor2_4 _3929_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1419_),
    .B(net20),
    .Y(_1673_));
 sky130_as_sc_hs__mux2_2 _3930_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1673_),
    .B(_1639_),
    .A(uio_out[0]),
    .Y(_1674_));
 sky130_as_sc_hs__buff_2 _3931_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1674_),
    .Y(_0267_));
 sky130_as_sc_hs__mux2_2 _3932_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1673_),
    .B(_1642_),
    .A(uio_out[1]),
    .Y(_1675_));
 sky130_as_sc_hs__buff_2 _3933_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1675_),
    .Y(_0268_));
 sky130_as_sc_hs__mux2_2 _3934_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1673_),
    .B(_1644_),
    .A(uio_out[2]),
    .Y(_1676_));
 sky130_as_sc_hs__buff_2 _3935_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1676_),
    .Y(_0269_));
 sky130_as_sc_hs__mux2_2 _3936_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1673_),
    .B(_1646_),
    .A(uio_out[3]),
    .Y(_1677_));
 sky130_as_sc_hs__buff_2 _3937_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1677_),
    .Y(_0270_));
 sky130_as_sc_hs__mux2_2 _3938_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1673_),
    .B(_1648_),
    .A(uio_out[4]),
    .Y(_1678_));
 sky130_as_sc_hs__buff_2 _3939_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1678_),
    .Y(_0271_));
 sky130_as_sc_hs__mux2_2 _3940_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1673_),
    .B(_1650_),
    .A(uio_out[5]),
    .Y(_1679_));
 sky130_as_sc_hs__buff_2 _3941_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1679_),
    .Y(_0272_));
 sky130_as_sc_hs__nor2_4 _3942_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1428_),
    .B(_1490_),
    .Y(_1680_));
 sky130_as_sc_hs__mux2_2 _3943_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1680_),
    .B(_1639_),
    .A(net331),
    .Y(_1681_));
 sky130_as_sc_hs__buff_2 _3944_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1681_),
    .Y(_0273_));
 sky130_as_sc_hs__mux2_2 _3945_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1680_),
    .B(_1642_),
    .A(net405),
    .Y(_1682_));
 sky130_as_sc_hs__buff_2 _3946_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1682_),
    .Y(_0274_));
 sky130_as_sc_hs__mux2_2 _3947_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1680_),
    .B(_1644_),
    .A(net512),
    .Y(_1683_));
 sky130_as_sc_hs__buff_2 _3948_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1683_),
    .Y(_0275_));
 sky130_as_sc_hs__mux2_2 _3949_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1680_),
    .B(_1646_),
    .A(net441),
    .Y(_1684_));
 sky130_as_sc_hs__buff_2 _3950_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1684_),
    .Y(_0276_));
 sky130_as_sc_hs__mux2_2 _3951_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1680_),
    .B(_1648_),
    .A(net446),
    .Y(_1685_));
 sky130_as_sc_hs__buff_2 _3952_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1685_),
    .Y(_0277_));
 sky130_as_sc_hs__mux2_2 _3953_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1680_),
    .B(_1650_),
    .A(net576),
    .Y(_1686_));
 sky130_as_sc_hs__buff_2 _3954_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1686_),
    .Y(_0278_));
 sky130_as_sc_hs__nor2_4 _3955_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1266_),
    .B(_1428_),
    .Y(_1687_));
 sky130_as_sc_hs__mux2_2 _3956_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1687_),
    .B(_1639_),
    .A(net349),
    .Y(_1688_));
 sky130_as_sc_hs__buff_2 _3957_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1688_),
    .Y(_0279_));
 sky130_as_sc_hs__mux2_2 _3958_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1687_),
    .B(_1642_),
    .A(net276),
    .Y(_1689_));
 sky130_as_sc_hs__buff_2 _3959_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1689_),
    .Y(_0280_));
 sky130_as_sc_hs__mux2_2 _3960_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1687_),
    .B(_1644_),
    .A(net408),
    .Y(_1690_));
 sky130_as_sc_hs__buff_2 _3961_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1690_),
    .Y(_0281_));
 sky130_as_sc_hs__mux2_2 _3962_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1687_),
    .B(_1646_),
    .A(net265),
    .Y(_1691_));
 sky130_as_sc_hs__buff_2 _3963_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1691_),
    .Y(_0282_));
 sky130_as_sc_hs__mux2_2 _3964_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1687_),
    .B(_1648_),
    .A(net418),
    .Y(_1692_));
 sky130_as_sc_hs__buff_2 _3965_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1692_),
    .Y(_0283_));
 sky130_as_sc_hs__mux2_2 _3966_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1687_),
    .B(_1650_),
    .A(net482),
    .Y(_1693_));
 sky130_as_sc_hs__buff_2 _3967_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1693_),
    .Y(_0284_));
 sky130_as_sc_hs__clkbuff_4 _3968_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1218_),
    .Y(_1694_));
 sky130_as_sc_hs__nor2_4 _3969_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1223_),
    .B(_1387_),
    .Y(_1695_));
 sky130_as_sc_hs__mux2_2 _3970_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1695_),
    .B(_1694_),
    .A(net339),
    .Y(_1696_));
 sky130_as_sc_hs__buff_2 _3971_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1696_),
    .Y(_0285_));
 sky130_as_sc_hs__clkbuff_4 _3972_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1230_),
    .Y(_1697_));
 sky130_as_sc_hs__mux2_2 _3973_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1695_),
    .B(_1697_),
    .A(net236),
    .Y(_1698_));
 sky130_as_sc_hs__buff_2 _3974_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1698_),
    .Y(_0286_));
 sky130_as_sc_hs__buff_4 _3975_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1235_),
    .Y(_1699_));
 sky130_as_sc_hs__mux2_2 _3976_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1695_),
    .B(_1699_),
    .A(net301),
    .Y(_1700_));
 sky130_as_sc_hs__buff_2 _3977_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1700_),
    .Y(_0287_));
 sky130_as_sc_hs__clkbuff_4 _3978_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1240_),
    .Y(_1701_));
 sky130_as_sc_hs__mux2_2 _3979_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1695_),
    .B(_1701_),
    .A(net403),
    .Y(_1702_));
 sky130_as_sc_hs__buff_2 _3980_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1702_),
    .Y(_0288_));
 sky130_as_sc_hs__buff_4 _3981_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1247_),
    .Y(_1703_));
 sky130_as_sc_hs__mux2_2 _3982_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1695_),
    .B(_1703_),
    .A(net583),
    .Y(_1704_));
 sky130_as_sc_hs__buff_2 _3983_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1704_),
    .Y(_0289_));
 sky130_as_sc_hs__buff_4 _3984_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1252_),
    .Y(_1705_));
 sky130_as_sc_hs__mux2_2 _3985_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1695_),
    .B(_1705_),
    .A(net386),
    .Y(_1706_));
 sky130_as_sc_hs__buff_2 _3986_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1706_),
    .Y(_0290_));
 sky130_as_sc_hs__nor2_4 _3987_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1427_),
    .B(net19),
    .Y(_1707_));
 sky130_as_sc_hs__mux2_2 _3988_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1707_),
    .B(_1694_),
    .A(net549),
    .Y(_1708_));
 sky130_as_sc_hs__buff_2 _3989_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1708_),
    .Y(_0291_));
 sky130_as_sc_hs__mux2_2 _3990_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1707_),
    .B(_1697_),
    .A(net467),
    .Y(_1709_));
 sky130_as_sc_hs__buff_2 _3991_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1709_),
    .Y(_0292_));
 sky130_as_sc_hs__mux2_2 _3992_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1707_),
    .B(_1699_),
    .A(net342),
    .Y(_1710_));
 sky130_as_sc_hs__buff_2 _3993_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1710_),
    .Y(_0293_));
 sky130_as_sc_hs__mux2_2 _3994_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1707_),
    .B(_1701_),
    .A(net531),
    .Y(_1711_));
 sky130_as_sc_hs__buff_2 _3995_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1711_),
    .Y(_0294_));
 sky130_as_sc_hs__mux2_2 _3996_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1707_),
    .B(_1703_),
    .A(net520),
    .Y(_1712_));
 sky130_as_sc_hs__buff_2 _3997_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1712_),
    .Y(_0295_));
 sky130_as_sc_hs__mux2_2 _3998_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1707_),
    .B(_1705_),
    .A(net240),
    .Y(_1713_));
 sky130_as_sc_hs__buff_2 _3999_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1713_),
    .Y(_0296_));
 sky130_as_sc_hs__nor2_4 _4000_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1366_),
    .B(_1387_),
    .Y(_1714_));
 sky130_as_sc_hs__mux2_2 _4001_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1714_),
    .B(_1694_),
    .A(net228),
    .Y(_1715_));
 sky130_as_sc_hs__buff_2 _4002_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1715_),
    .Y(_0297_));
 sky130_as_sc_hs__mux2_2 _4003_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1714_),
    .B(_1697_),
    .A(net284),
    .Y(_1716_));
 sky130_as_sc_hs__buff_2 _4004_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1716_),
    .Y(_0298_));
 sky130_as_sc_hs__mux2_2 _4005_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1714_),
    .B(_1699_),
    .A(net320),
    .Y(_1717_));
 sky130_as_sc_hs__buff_2 _4006_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1717_),
    .Y(_0299_));
 sky130_as_sc_hs__mux2_2 _4007_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1714_),
    .B(_1701_),
    .A(net377),
    .Y(_1718_));
 sky130_as_sc_hs__buff_2 _4008_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1718_),
    .Y(_0300_));
 sky130_as_sc_hs__mux2_2 _4009_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1714_),
    .B(_1703_),
    .A(net231),
    .Y(_1719_));
 sky130_as_sc_hs__buff_2 _4010_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1719_),
    .Y(_0301_));
 sky130_as_sc_hs__mux2_2 _4011_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1714_),
    .B(_1705_),
    .A(net410),
    .Y(_1720_));
 sky130_as_sc_hs__buff_2 _4012_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1720_),
    .Y(_0302_));
 sky130_as_sc_hs__nor2_4 _4013_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1402_),
    .B(_1554_),
    .Y(_1721_));
 sky130_as_sc_hs__mux2_2 _4014_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1721_),
    .B(_1694_),
    .A(net572),
    .Y(_1722_));
 sky130_as_sc_hs__buff_2 _4015_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1722_),
    .Y(_0303_));
 sky130_as_sc_hs__mux2_2 _4016_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1721_),
    .B(_1697_),
    .A(net371),
    .Y(_1723_));
 sky130_as_sc_hs__buff_2 _4017_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1723_),
    .Y(_0304_));
 sky130_as_sc_hs__mux2_2 _4018_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1721_),
    .B(_1699_),
    .A(net480),
    .Y(_1724_));
 sky130_as_sc_hs__buff_2 _4019_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1724_),
    .Y(_0305_));
 sky130_as_sc_hs__mux2_2 _4020_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1721_),
    .B(_1701_),
    .A(net370),
    .Y(_1725_));
 sky130_as_sc_hs__buff_2 _4021_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1725_),
    .Y(_0306_));
 sky130_as_sc_hs__mux2_2 _4022_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1721_),
    .B(_1703_),
    .A(net456),
    .Y(_1726_));
 sky130_as_sc_hs__buff_2 _4023_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1726_),
    .Y(_0307_));
 sky130_as_sc_hs__mux2_2 _4024_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1721_),
    .B(_1705_),
    .A(net523),
    .Y(_1727_));
 sky130_as_sc_hs__buff_2 _4025_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1727_),
    .Y(_0308_));
 sky130_as_sc_hs__nor2_4 _4026_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1387_),
    .B(_1490_),
    .Y(_1728_));
 sky130_as_sc_hs__mux2_2 _4027_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1728_),
    .B(_1694_),
    .A(net264),
    .Y(_1729_));
 sky130_as_sc_hs__buff_2 _4028_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1729_),
    .Y(_0309_));
 sky130_as_sc_hs__mux2_2 _4029_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1728_),
    .B(_1697_),
    .A(net409),
    .Y(_1730_));
 sky130_as_sc_hs__buff_2 _4030_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1730_),
    .Y(_0310_));
 sky130_as_sc_hs__mux2_2 _4031_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1728_),
    .B(_1699_),
    .A(net542),
    .Y(_1731_));
 sky130_as_sc_hs__buff_2 _4032_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1731_),
    .Y(_0311_));
 sky130_as_sc_hs__mux2_2 _4033_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1728_),
    .B(_1701_),
    .A(net268),
    .Y(_1732_));
 sky130_as_sc_hs__buff_2 _4034_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1732_),
    .Y(_0312_));
 sky130_as_sc_hs__mux2_2 _4035_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1728_),
    .B(_1703_),
    .A(net429),
    .Y(_1733_));
 sky130_as_sc_hs__buff_2 _4036_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1733_),
    .Y(_0313_));
 sky130_as_sc_hs__mux2_2 _4037_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1728_),
    .B(_1705_),
    .A(net346),
    .Y(_1734_));
 sky130_as_sc_hs__buff_2 _4038_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1734_),
    .Y(_0314_));
 sky130_as_sc_hs__clkbuff_4 _4039_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1156_),
    .Y(_1735_));
 sky130_as_sc_hs__aoi21_2 _4040_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0607_),
    .B(net21),
    .C(_1130_),
    .Y(_1736_));
 sky130_as_sc_hs__nor2_4 _4041_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1365_),
    .B(net18),
    .Y(_1737_));
 sky130_as_sc_hs__mux2_2 _4042_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1737_),
    .B(_1217_),
    .A(uio_oe[0]),
    .Y(_1738_));
 sky130_as_sc_hs__or2_2 _4043_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1735_),
    .B(_1738_),
    .Y(_1739_));
 sky130_as_sc_hs__buff_2 _4044_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1739_),
    .Y(_0315_));
 sky130_as_sc_hs__mux2_2 _4045_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1737_),
    .B(_1229_),
    .A(uio_oe[1]),
    .Y(_1740_));
 sky130_as_sc_hs__or2_2 _4046_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1735_),
    .B(_1740_),
    .Y(_1741_));
 sky130_as_sc_hs__buff_2 _4047_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1741_),
    .Y(_0316_));
 sky130_as_sc_hs__mux2_2 _4048_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1737_),
    .B(_1234_),
    .A(uio_oe[2]),
    .Y(_1742_));
 sky130_as_sc_hs__or2_2 _4049_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1735_),
    .B(_1742_),
    .Y(_1743_));
 sky130_as_sc_hs__buff_2 _4050_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1743_),
    .Y(_0317_));
 sky130_as_sc_hs__mux2_2 _4051_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1737_),
    .B(_1239_),
    .A(uio_oe[3]),
    .Y(_1744_));
 sky130_as_sc_hs__or2_2 _4052_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1157_),
    .B(_1744_),
    .Y(_1745_));
 sky130_as_sc_hs__buff_2 _4053_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1745_),
    .Y(_0318_));
 sky130_as_sc_hs__mux2_2 _4054_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1737_),
    .B(_1246_),
    .A(uio_oe[4]),
    .Y(_1746_));
 sky130_as_sc_hs__or2_2 _4055_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1157_),
    .B(_1746_),
    .Y(_1747_));
 sky130_as_sc_hs__buff_2 _4056_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1747_),
    .Y(_0319_));
 sky130_as_sc_hs__mux2_2 _4057_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1737_),
    .B(_1251_),
    .A(uio_oe[5]),
    .Y(_1748_));
 sky130_as_sc_hs__or2_2 _4058_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1157_),
    .B(_1748_),
    .Y(_1749_));
 sky130_as_sc_hs__buff_2 _4059_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1749_),
    .Y(_0320_));
 sky130_as_sc_hs__nor2_4 _4060_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1402_),
    .B(_1428_),
    .Y(_1750_));
 sky130_as_sc_hs__mux2_2 _4061_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1750_),
    .B(_1694_),
    .A(net477),
    .Y(_1751_));
 sky130_as_sc_hs__buff_2 _4062_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1751_),
    .Y(_0321_));
 sky130_as_sc_hs__mux2_2 _4063_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1750_),
    .B(_1697_),
    .A(net217),
    .Y(_1752_));
 sky130_as_sc_hs__buff_2 _4064_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1752_),
    .Y(_0322_));
 sky130_as_sc_hs__mux2_2 _4065_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1750_),
    .B(_1699_),
    .A(net398),
    .Y(_1753_));
 sky130_as_sc_hs__buff_2 _4066_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1753_),
    .Y(_0323_));
 sky130_as_sc_hs__mux2_2 _4067_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1750_),
    .B(_1701_),
    .A(net391),
    .Y(_1754_));
 sky130_as_sc_hs__buff_2 _4068_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1754_),
    .Y(_0324_));
 sky130_as_sc_hs__mux2_2 _4069_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1750_),
    .B(_1703_),
    .A(net457),
    .Y(_1755_));
 sky130_as_sc_hs__buff_2 _4070_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1755_),
    .Y(_0325_));
 sky130_as_sc_hs__mux2_2 _4071_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1750_),
    .B(_1705_),
    .A(net437),
    .Y(_1756_));
 sky130_as_sc_hs__buff_2 _4072_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1756_),
    .Y(_0326_));
 sky130_as_sc_hs__nor2_4 _4073_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1275_),
    .B(_1387_),
    .Y(_1757_));
 sky130_as_sc_hs__mux2_2 _4074_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1757_),
    .B(_1694_),
    .A(net310),
    .Y(_1758_));
 sky130_as_sc_hs__buff_2 _4075_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1758_),
    .Y(_0327_));
 sky130_as_sc_hs__mux2_2 _4076_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1757_),
    .B(_1697_),
    .A(net271),
    .Y(_1759_));
 sky130_as_sc_hs__buff_2 _4077_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1759_),
    .Y(_0328_));
 sky130_as_sc_hs__mux2_2 _4078_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1757_),
    .B(_1699_),
    .A(net368),
    .Y(_1760_));
 sky130_as_sc_hs__buff_2 _4079_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1760_),
    .Y(_0329_));
 sky130_as_sc_hs__mux2_2 _4080_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1757_),
    .B(_1701_),
    .A(net483),
    .Y(_1761_));
 sky130_as_sc_hs__buff_2 _4081_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1761_),
    .Y(_0330_));
 sky130_as_sc_hs__mux2_2 _4082_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1757_),
    .B(_1703_),
    .A(net401),
    .Y(_1762_));
 sky130_as_sc_hs__buff_2 _4083_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1762_),
    .Y(_0331_));
 sky130_as_sc_hs__mux2_2 _4084_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1757_),
    .B(_1705_),
    .A(net202),
    .Y(_1763_));
 sky130_as_sc_hs__buff_2 _4085_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1763_),
    .Y(_0332_));
 sky130_as_sc_hs__nor2_4 _4086_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1222_),
    .B(net18),
    .Y(_1764_));
 sky130_as_sc_hs__mux2_2 _4087_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1764_),
    .B(_1470_),
    .A(uo_out[0]),
    .Y(_1765_));
 sky130_as_sc_hs__and2_2 _4088_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net147),
    .B(_1765_),
    .Y(_1766_));
 sky130_as_sc_hs__buff_2 _4089_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1766_),
    .Y(_0333_));
 sky130_as_sc_hs__mux2_2 _4090_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1764_),
    .B(_1475_),
    .A(uo_out[1]),
    .Y(_1767_));
 sky130_as_sc_hs__and2_2 _4091_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net147),
    .B(_1767_),
    .Y(_1768_));
 sky130_as_sc_hs__buff_2 _4092_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1768_),
    .Y(_0334_));
 sky130_as_sc_hs__mux2_2 _4093_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1764_),
    .B(_1478_),
    .A(uo_out[2]),
    .Y(_1769_));
 sky130_as_sc_hs__and2_2 _4094_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net147),
    .B(_1769_),
    .Y(_1770_));
 sky130_as_sc_hs__buff_2 _4095_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1770_),
    .Y(_0335_));
 sky130_as_sc_hs__mux2_2 _4096_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1764_),
    .B(_1481_),
    .A(uo_out[3]),
    .Y(_1771_));
 sky130_as_sc_hs__and2_2 _4097_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net147),
    .B(_1771_),
    .Y(_1772_));
 sky130_as_sc_hs__buff_2 _4098_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1772_),
    .Y(_0336_));
 sky130_as_sc_hs__mux2_2 _4099_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1764_),
    .B(_1484_),
    .A(uo_out[4]),
    .Y(_1773_));
 sky130_as_sc_hs__and2_2 _4100_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net147),
    .B(_1773_),
    .Y(_1774_));
 sky130_as_sc_hs__buff_2 _4101_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1774_),
    .Y(_0337_));
 sky130_as_sc_hs__mux2_2 _4102_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1764_),
    .B(_1487_),
    .A(uo_out[5]),
    .Y(_1775_));
 sky130_as_sc_hs__and2_2 _4103_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net147),
    .B(_1775_),
    .Y(_1776_));
 sky130_as_sc_hs__buff_2 _4104_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1776_),
    .Y(_0338_));
 sky130_as_sc_hs__clkbuff_4 _4105_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1217_),
    .Y(_1777_));
 sky130_as_sc_hs__nor2_4 _4106_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1490_),
    .B(_1554_),
    .Y(_1778_));
 sky130_as_sc_hs__mux2_2 _4107_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1778_),
    .B(_1777_),
    .A(net209),
    .Y(_1779_));
 sky130_as_sc_hs__buff_2 _4108_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1779_),
    .Y(_0339_));
 sky130_as_sc_hs__buff_4 _4109_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1229_),
    .Y(_1780_));
 sky130_as_sc_hs__mux2_2 _4110_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1778_),
    .B(_1780_),
    .A(net385),
    .Y(_1781_));
 sky130_as_sc_hs__buff_2 _4111_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1781_),
    .Y(_0340_));
 sky130_as_sc_hs__buff_4 _4112_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1234_),
    .Y(_1782_));
 sky130_as_sc_hs__mux2_2 _4113_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1778_),
    .B(_1782_),
    .A(net258),
    .Y(_1783_));
 sky130_as_sc_hs__buff_2 _4114_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1783_),
    .Y(_0341_));
 sky130_as_sc_hs__clkbuff_4 _4115_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1239_),
    .Y(_1784_));
 sky130_as_sc_hs__mux2_2 _4116_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1778_),
    .B(_1784_),
    .A(net463),
    .Y(_1785_));
 sky130_as_sc_hs__buff_2 _4117_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1785_),
    .Y(_0342_));
 sky130_as_sc_hs__clkbuff_4 _4118_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1246_),
    .Y(_1786_));
 sky130_as_sc_hs__mux2_2 _4119_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1778_),
    .B(_1786_),
    .A(net396),
    .Y(_1787_));
 sky130_as_sc_hs__buff_2 _4120_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1787_),
    .Y(_0343_));
 sky130_as_sc_hs__buff_4 _4121_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1251_),
    .Y(_1788_));
 sky130_as_sc_hs__mux2_2 _4122_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1778_),
    .B(_1788_),
    .A(net372),
    .Y(_1789_));
 sky130_as_sc_hs__buff_2 _4123_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1789_),
    .Y(_0344_));
 sky130_as_sc_hs__nor2_4 _4124_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1401_),
    .B(_1736_),
    .Y(_1790_));
 sky130_as_sc_hs__mux2_2 _4125_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1790_),
    .B(_1777_),
    .A(net532),
    .Y(_1791_));
 sky130_as_sc_hs__buff_2 _4126_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1791_),
    .Y(_0345_));
 sky130_as_sc_hs__mux2_2 _4127_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1790_),
    .B(_1780_),
    .A(net204),
    .Y(_1792_));
 sky130_as_sc_hs__buff_2 _4128_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1792_),
    .Y(_0346_));
 sky130_as_sc_hs__mux2_2 _4129_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1790_),
    .B(_1782_),
    .A(net528),
    .Y(_1793_));
 sky130_as_sc_hs__buff_2 _4130_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1793_),
    .Y(_0347_));
 sky130_as_sc_hs__mux2_2 _4131_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1790_),
    .B(_1784_),
    .A(net199),
    .Y(_1794_));
 sky130_as_sc_hs__buff_2 _4132_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1794_),
    .Y(_0348_));
 sky130_as_sc_hs__mux2_2 _4133_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1790_),
    .B(_1786_),
    .A(net433),
    .Y(_1795_));
 sky130_as_sc_hs__buff_2 _4134_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1795_),
    .Y(_0349_));
 sky130_as_sc_hs__mux2_2 _4135_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1790_),
    .B(_1788_),
    .A(net402),
    .Y(_1796_));
 sky130_as_sc_hs__buff_2 _4136_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1796_),
    .Y(_0350_));
 sky130_as_sc_hs__nor2_4 _4137_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1256_),
    .B(_1428_),
    .Y(_1797_));
 sky130_as_sc_hs__mux2_2 _4138_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1797_),
    .B(_1777_),
    .A(net473),
    .Y(_1798_));
 sky130_as_sc_hs__buff_2 _4139_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1798_),
    .Y(_0351_));
 sky130_as_sc_hs__mux2_2 _4140_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1797_),
    .B(_1780_),
    .A(net393),
    .Y(_1799_));
 sky130_as_sc_hs__buff_2 _4141_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1799_),
    .Y(_0352_));
 sky130_as_sc_hs__mux2_2 _4142_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1797_),
    .B(_1782_),
    .A(net270),
    .Y(_1800_));
 sky130_as_sc_hs__buff_2 _4143_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1800_),
    .Y(_0353_));
 sky130_as_sc_hs__mux2_2 _4144_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1797_),
    .B(_1784_),
    .A(net492),
    .Y(_1801_));
 sky130_as_sc_hs__buff_2 _4145_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1801_),
    .Y(_0354_));
 sky130_as_sc_hs__mux2_2 _4146_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1797_),
    .B(_1786_),
    .A(net502),
    .Y(_1802_));
 sky130_as_sc_hs__buff_2 _4147_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1802_),
    .Y(_0355_));
 sky130_as_sc_hs__mux2_2 _4148_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1797_),
    .B(_1788_),
    .A(net543),
    .Y(_1803_));
 sky130_as_sc_hs__buff_2 _4149_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1803_),
    .Y(_0356_));
 sky130_as_sc_hs__nor2_4 _4150_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1386_),
    .B(_1402_),
    .Y(_1804_));
 sky130_as_sc_hs__mux2_2 _4151_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1804_),
    .B(_1777_),
    .A(net253),
    .Y(_1805_));
 sky130_as_sc_hs__buff_2 _4152_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1805_),
    .Y(_0357_));
 sky130_as_sc_hs__mux2_2 _4153_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1804_),
    .B(_1780_),
    .A(net431),
    .Y(_1806_));
 sky130_as_sc_hs__buff_2 _4154_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1806_),
    .Y(_0358_));
 sky130_as_sc_hs__mux2_2 _4155_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1804_),
    .B(_1782_),
    .A(net454),
    .Y(_1807_));
 sky130_as_sc_hs__buff_2 _4156_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1807_),
    .Y(_0359_));
 sky130_as_sc_hs__mux2_2 _4157_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1804_),
    .B(_1784_),
    .A(net343),
    .Y(_1808_));
 sky130_as_sc_hs__buff_2 _4158_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1808_),
    .Y(_0360_));
 sky130_as_sc_hs__mux2_2 _4159_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1804_),
    .B(_1786_),
    .A(net412),
    .Y(_1809_));
 sky130_as_sc_hs__buff_2 _4160_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1809_),
    .Y(_0361_));
 sky130_as_sc_hs__mux2_2 _4161_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1804_),
    .B(_1788_),
    .A(net425),
    .Y(_1810_));
 sky130_as_sc_hs__buff_2 _4162_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1810_),
    .Y(_0362_));
 sky130_as_sc_hs__nor2_4 _4163_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1366_),
    .B(_1554_),
    .Y(_1811_));
 sky130_as_sc_hs__mux2_2 _4164_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1811_),
    .B(_1777_),
    .A(net280),
    .Y(_1812_));
 sky130_as_sc_hs__buff_2 _4165_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1812_),
    .Y(_0363_));
 sky130_as_sc_hs__mux2_2 _4166_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1811_),
    .B(_1780_),
    .A(net503),
    .Y(_1813_));
 sky130_as_sc_hs__buff_2 _4167_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1813_),
    .Y(_0364_));
 sky130_as_sc_hs__mux2_2 _4168_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1811_),
    .B(_1782_),
    .A(net324),
    .Y(_1814_));
 sky130_as_sc_hs__buff_2 _4169_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1814_),
    .Y(_0365_));
 sky130_as_sc_hs__mux2_2 _4170_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1811_),
    .B(_1784_),
    .A(net279),
    .Y(_1815_));
 sky130_as_sc_hs__buff_2 _4171_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1815_),
    .Y(_0366_));
 sky130_as_sc_hs__mux2_2 _4172_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1811_),
    .B(_1786_),
    .A(net249),
    .Y(_1816_));
 sky130_as_sc_hs__buff_2 _4173_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1816_),
    .Y(_0367_));
 sky130_as_sc_hs__mux2_2 _4174_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1811_),
    .B(_1788_),
    .A(net550),
    .Y(_1817_));
 sky130_as_sc_hs__buff_2 _4175_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1817_),
    .Y(_0368_));
 sky130_as_sc_hs__nor2_4 _4176_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1368_),
    .B(net19),
    .Y(_1818_));
 sky130_as_sc_hs__mux2_2 _4177_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1818_),
    .B(_1777_),
    .A(net200),
    .Y(_1819_));
 sky130_as_sc_hs__buff_2 _4178_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1819_),
    .Y(_0369_));
 sky130_as_sc_hs__mux2_2 _4179_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1818_),
    .B(_1780_),
    .A(net493),
    .Y(_1820_));
 sky130_as_sc_hs__buff_2 _4180_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1820_),
    .Y(_0370_));
 sky130_as_sc_hs__mux2_2 _4181_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1818_),
    .B(_1782_),
    .A(net544),
    .Y(_1821_));
 sky130_as_sc_hs__buff_2 _4182_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1821_),
    .Y(_0371_));
 sky130_as_sc_hs__mux2_2 _4183_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1818_),
    .B(_1784_),
    .A(net435),
    .Y(_1822_));
 sky130_as_sc_hs__buff_2 _4184_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1822_),
    .Y(_0372_));
 sky130_as_sc_hs__mux2_2 _4185_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1818_),
    .B(_1786_),
    .A(net588),
    .Y(_1823_));
 sky130_as_sc_hs__buff_2 _4186_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1823_),
    .Y(_0373_));
 sky130_as_sc_hs__mux2_2 _4187_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1818_),
    .B(_1788_),
    .A(net334),
    .Y(_1824_));
 sky130_as_sc_hs__buff_2 _4188_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1824_),
    .Y(_0374_));
 sky130_as_sc_hs__nor2_4 _4189_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1223_),
    .B(_1554_),
    .Y(_1825_));
 sky130_as_sc_hs__mux2_2 _4190_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1825_),
    .B(_1777_),
    .A(net430),
    .Y(_1826_));
 sky130_as_sc_hs__buff_2 _4191_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1826_),
    .Y(_0375_));
 sky130_as_sc_hs__mux2_2 _4192_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1825_),
    .B(_1780_),
    .A(net267),
    .Y(_1827_));
 sky130_as_sc_hs__buff_2 _4193_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1827_),
    .Y(_0376_));
 sky130_as_sc_hs__mux2_2 _4194_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1825_),
    .B(_1782_),
    .A(net384),
    .Y(_1828_));
 sky130_as_sc_hs__buff_2 _4195_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1828_),
    .Y(_0377_));
 sky130_as_sc_hs__mux2_2 _4196_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1825_),
    .B(_1784_),
    .A(net238),
    .Y(_1829_));
 sky130_as_sc_hs__buff_2 _4197_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1829_),
    .Y(_0378_));
 sky130_as_sc_hs__mux2_2 _4198_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1825_),
    .B(_1786_),
    .A(net272),
    .Y(_1830_));
 sky130_as_sc_hs__buff_2 _4199_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1830_),
    .Y(_0379_));
 sky130_as_sc_hs__mux2_2 _4200_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1825_),
    .B(_1788_),
    .A(net315),
    .Y(_1831_));
 sky130_as_sc_hs__buff_2 _4201_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1831_),
    .Y(_0380_));
 sky130_as_sc_hs__nor2_4 _4202_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1265_),
    .B(_1369_),
    .Y(_1832_));
 sky130_as_sc_hs__mux2_2 _4203_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1832_),
    .B(_1470_),
    .A(net462),
    .Y(_1833_));
 sky130_as_sc_hs__buff_2 _4204_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1833_),
    .Y(_0381_));
 sky130_as_sc_hs__mux2_2 _4205_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1832_),
    .B(_1475_),
    .A(net214),
    .Y(_1834_));
 sky130_as_sc_hs__buff_2 _4206_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1834_),
    .Y(_0382_));
 sky130_as_sc_hs__mux2_2 _4207_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1832_),
    .B(_1478_),
    .A(net400),
    .Y(_1835_));
 sky130_as_sc_hs__buff_2 _4208_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1835_),
    .Y(_0383_));
 sky130_as_sc_hs__mux2_2 _4209_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1832_),
    .B(_1481_),
    .A(net188),
    .Y(_1836_));
 sky130_as_sc_hs__buff_2 _4210_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1836_),
    .Y(_0384_));
 sky130_as_sc_hs__mux2_2 _4211_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1832_),
    .B(_1484_),
    .A(net469),
    .Y(_1837_));
 sky130_as_sc_hs__buff_2 _4212_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1837_),
    .Y(_0385_));
 sky130_as_sc_hs__mux2_2 _4213_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1832_),
    .B(_1487_),
    .A(net395),
    .Y(_1838_));
 sky130_as_sc_hs__buff_2 _4214_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1838_),
    .Y(_0386_));
 sky130_as_sc_hs__nor2_4 _4215_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1256_),
    .B(_1554_),
    .Y(_1839_));
 sky130_as_sc_hs__mux2_2 _4216_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1839_),
    .B(_1470_),
    .A(net415),
    .Y(_1840_));
 sky130_as_sc_hs__buff_2 _4217_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1840_),
    .Y(_0387_));
 sky130_as_sc_hs__mux2_2 _4218_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1839_),
    .B(_1475_),
    .A(net445),
    .Y(_1841_));
 sky130_as_sc_hs__buff_2 _4219_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1841_),
    .Y(_0388_));
 sky130_as_sc_hs__mux2_2 _4220_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1839_),
    .B(_1478_),
    .A(net222),
    .Y(_1842_));
 sky130_as_sc_hs__buff_2 _4221_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1842_),
    .Y(_0389_));
 sky130_as_sc_hs__mux2_2 _4222_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1839_),
    .B(_1481_),
    .A(net413),
    .Y(_1843_));
 sky130_as_sc_hs__buff_2 _4223_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1843_),
    .Y(_0390_));
 sky130_as_sc_hs__mux2_2 _4224_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1839_),
    .B(_1484_),
    .A(net347),
    .Y(_1844_));
 sky130_as_sc_hs__buff_2 _4225_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1844_),
    .Y(_0391_));
 sky130_as_sc_hs__mux2_2 _4226_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1839_),
    .B(_1487_),
    .A(net491),
    .Y(_1845_));
 sky130_as_sc_hs__buff_2 _4227_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1845_),
    .Y(_0392_));
 sky130_as_sc_hs__nor2_4 _4228_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1255_),
    .B(net18),
    .Y(_1846_));
 sky130_as_sc_hs__mux2_2 _4229_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1846_),
    .B(_1470_),
    .A(net416),
    .Y(_1847_));
 sky130_as_sc_hs__buff_2 _4230_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1847_),
    .Y(_0393_));
 sky130_as_sc_hs__mux2_2 _4231_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1846_),
    .B(_1475_),
    .A(net250),
    .Y(_1848_));
 sky130_as_sc_hs__buff_2 _4232_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1848_),
    .Y(_0394_));
 sky130_as_sc_hs__mux2_2 _4233_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1846_),
    .B(_1478_),
    .A(net452),
    .Y(_1849_));
 sky130_as_sc_hs__buff_2 _4234_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1849_),
    .Y(_0395_));
 sky130_as_sc_hs__mux2_2 _4235_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1846_),
    .B(_1481_),
    .A(net244),
    .Y(_1850_));
 sky130_as_sc_hs__buff_2 _4236_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1850_),
    .Y(_0396_));
 sky130_as_sc_hs__mux2_2 _4237_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1846_),
    .B(_1484_),
    .A(net421),
    .Y(_1851_));
 sky130_as_sc_hs__buff_2 _4238_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1851_),
    .Y(_0397_));
 sky130_as_sc_hs__mux2_2 _4239_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1846_),
    .B(_1487_),
    .A(net375),
    .Y(_1852_));
 sky130_as_sc_hs__buff_2 _4240_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1852_),
    .Y(_0398_));
 sky130_as_sc_hs__ao21_2 _4241_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0679_),
    .B(_0947_),
    .C(_0958_),
    .Y(_1853_));
 sky130_as_sc_hs__nor2_2 _4242_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0936_),
    .B(_0943_),
    .Y(_1854_));
 sky130_as_sc_hs__iao211_2 _4243_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1853_),
    .B(_0951_),
    .C(_0928_),
    .D(_1854_),
    .Y(_1855_));
 sky130_as_sc_hs__nand2_2 _4244_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net23),
    .B(_0927_),
    .Y(_1856_));
 sky130_as_sc_hs__nand2_2 _4245_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0967_),
    .B(_0975_),
    .Y(_1857_));
 sky130_as_sc_hs__nand4_2 _4246_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net23),
    .B(_0927_),
    .C(_0985_),
    .Y(_1858_),
    .D(_0995_));
 sky130_as_sc_hs__oa22_2 _4247_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1856_),
    .B(_0960_),
    .C(_1857_),
    .D(_1858_),
    .Y(_1859_));
 sky130_as_sc_hs__inv_2 _4248_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_0998_),
    .Y(_1860_));
 sky130_as_sc_hs__inv_2 _4249_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net132),
    .Y(_1861_));
 sky130_as_sc_hs__aoi31_2 _4250_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1855_),
    .B(_1859_),
    .C(_1860_),
    .D(_1861_),
    .Y(_1862_));
 sky130_as_sc_hs__inv_2 _4251_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(carry),
    .Y(_1863_));
 sky130_as_sc_hs__nand2_2 _4252_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1863_),
    .B(net43),
    .Y(_1864_));
 sky130_as_sc_hs__inv_2 _4253_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_1864_),
    .Y(_1865_));
 sky130_as_sc_hs__aoi211_2 _4254_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_0997_),
    .C(_0998_),
    .D(net132),
    .Y(_1866_),
    .A(_0928_));
 sky130_as_sc_hs__nor2_2 _4255_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net17),
    .B(_1866_),
    .Y(_1867_));
 sky130_as_sc_hs__nand2_2 _4256_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(carry),
    .B(_1128_),
    .Y(_1868_));
 sky130_as_sc_hs__or2_2 _4257_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net133),
    .B(_1864_),
    .Y(_1869_));
 sky130_as_sc_hs__oai22_2 _4258_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1867_),
    .B(_1868_),
    .C(_1869_),
    .D(_0999_),
    .Y(_1870_));
 sky130_as_sc_hs__ao22_2 _4259_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net17),
    .C(_1870_),
    .B(_1865_),
    .D(net37),
    .Y(_1871_));
 sky130_as_sc_hs__ao31_2 _4260_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net37),
    .B(_1868_),
    .C(_1864_),
    .D(_1123_),
    .Y(_1872_));
 sky130_as_sc_hs__ao21_2 _4261_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1133_),
    .B(net17),
    .C(_1001_),
    .Y(_1873_));
 sky130_as_sc_hs__ao22_2 _4262_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1867_),
    .C(_1873_),
    .B(_1872_),
    .D(_1151_),
    .Y(_1874_));
 sky130_as_sc_hs__ao21_2 _4263_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net46),
    .B(_1871_),
    .C(_1874_),
    .Y(_1875_));
 sky130_as_sc_hs__xnor2_2 _4264_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net124),
    .Y(_1876_),
    .B(_0918_));
 sky130_as_sc_hs__and2_2 _4265_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net126),
    .B(_0840_),
    .Y(_1877_));
 sky130_as_sc_hs__nor2_2 _4266_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net127),
    .B(_0840_),
    .Y(_1878_));
 sky130_as_sc_hs__nor2_4 _4267_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1877_),
    .B(_1878_),
    .Y(_1879_));
 sky130_as_sc_hs__inv_2 _4268_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\A[3] ),
    .Y(_1880_));
 sky130_as_sc_hs__xnor2_2 _4269_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1880_),
    .Y(_1881_),
    .B(_0753_));
 sky130_as_sc_hs__xnor2_2 _4270_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net128),
    .Y(_1882_),
    .B(_0646_));
 sky130_as_sc_hs__aoi211_2 _4271_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1081_),
    .C(_1082_),
    .D(net130),
    .Y(_1883_),
    .A(_1016_));
 sky130_as_sc_hs__nand2_2 _4272_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1016_),
    .B(_1080_),
    .Y(_1884_));
 sky130_as_sc_hs__nand3_2 _4273_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1016_),
    .B(_1032_),
    .C(_1048_),
    .Y(_1885_));
 sky130_as_sc_hs__inv_2 _4274_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_1082_),
    .Y(_1886_));
 sky130_as_sc_hs__inv_2 _4275_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net131),
    .Y(_1887_));
 sky130_as_sc_hs__aoi31_2 _4276_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1884_),
    .B(_1885_),
    .C(_1886_),
    .D(_1887_),
    .Y(_1888_));
 sky130_as_sc_hs__oa22_2 _4277_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net17),
    .B(_1866_),
    .C(_1883_),
    .D(_1888_),
    .Y(_1889_));
 sky130_as_sc_hs__buff_2 _4278_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1889_),
    .Y(_1890_));
 sky130_as_sc_hs__nand3_2 _4279_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1881_),
    .B(_1882_),
    .C(_1890_),
    .Y(_1891_));
 sky130_as_sc_hs__inv_2 _4280_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_1891_),
    .Y(_1892_));
 sky130_as_sc_hs__nand3_2 _4281_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1151_),
    .B(_1182_),
    .C(_1129_),
    .Y(_1893_));
 sky130_as_sc_hs__ao31_2 _4282_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1876_),
    .B(_1879_),
    .C(_1892_),
    .D(_1893_),
    .Y(_1894_));
 sky130_as_sc_hs__nand2_2 _4283_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1150_),
    .B(net45),
    .Y(_1895_));
 sky130_as_sc_hs__nor2_2 _4284_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net41),
    .B(_1895_),
    .Y(_1896_));
 sky130_as_sc_hs__ao31_2 _4285_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net128),
    .B(_1093_),
    .C(_0753_),
    .D(\A[3] ),
    .Y(_1897_));
 sky130_as_sc_hs__ao21_2 _4286_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net128),
    .B(_1094_),
    .C(_0753_),
    .Y(_1898_));
 sky130_as_sc_hs__nand2_2 _4287_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1897_),
    .B(_1898_),
    .Y(_1899_));
 sky130_as_sc_hs__buff_2 _4288_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1899_),
    .Y(_1900_));
 sky130_as_sc_hs__aoi21_2 _4289_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1016_),
    .B(_1081_),
    .C(_1082_),
    .Y(_1901_));
 sky130_as_sc_hs__ao31_2 _4290_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1855_),
    .B(_1859_),
    .C(_1860_),
    .D(net132),
    .Y(_1902_));
 sky130_as_sc_hs__maj3_2 _4291_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1901_),
    .A(net130),
    .C(_1902_),
    .Y(_1903_));
 sky130_as_sc_hs__nand3_2 _4292_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1881_),
    .B(_1882_),
    .C(_1903_),
    .Y(_1904_));
 sky130_as_sc_hs__buff_2 _4293_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1904_),
    .Y(_1905_));
 sky130_as_sc_hs__clkbuff_4 _4294_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1882_),
    .Y(_1906_));
 sky130_as_sc_hs__buff_4 _4295_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0840_),
    .Y(_1907_));
 sky130_as_sc_hs__iao211_2 _4296_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0883_),
    .B(_0884_),
    .C(_0917_),
    .D(_1907_),
    .Y(_1908_));
 sky130_as_sc_hs__ao31_2 _4297_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1881_),
    .B(_1906_),
    .C(_1890_),
    .D(_1908_),
    .Y(_1909_));
 sky130_as_sc_hs__clkbuff_4 _4298_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1881_),
    .Y(_1910_));
 sky130_as_sc_hs__iao211_2 _4299_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0883_),
    .B(_0884_),
    .C(_0917_),
    .D(net126),
    .Y(_1911_));
 sky130_as_sc_hs__ao31_2 _4300_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1910_),
    .B(_1906_),
    .C(_1890_),
    .D(_1911_),
    .Y(_1912_));
 sky130_as_sc_hs__ao22_2 _4301_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1900_),
    .C(_1909_),
    .B(_1905_),
    .D(_1912_),
    .Y(_1913_));
 sky130_as_sc_hs__nand2_2 _4302_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net125),
    .B(_1907_),
    .Y(_1914_));
 sky130_as_sc_hs__ao31_2 _4303_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1910_),
    .B(_1906_),
    .C(_1890_),
    .D(_1914_),
    .Y(_1915_));
 sky130_as_sc_hs__nand2_2 _4304_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net124),
    .B(net127),
    .Y(_1916_));
 sky130_as_sc_hs__ao31_2 _4305_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1910_),
    .B(_1906_),
    .C(_1890_),
    .D(_1916_),
    .Y(_1917_));
 sky130_as_sc_hs__ao22_2 _4306_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1900_),
    .C(_1915_),
    .B(_1905_),
    .D(_1917_),
    .Y(_1918_));
 sky130_as_sc_hs__inv_2 _4307_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net125),
    .Y(_1919_));
 sky130_as_sc_hs__nand2_2 _4308_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net127),
    .B(_1907_),
    .Y(_1920_));
 sky130_as_sc_hs__ao21_2 _4309_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1919_),
    .B(_1920_),
    .C(_0918_),
    .Y(_1921_));
 sky130_as_sc_hs__oa21_2 _4310_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0842_),
    .B(_1916_),
    .C(_1921_),
    .Y(_1922_));
 sky130_as_sc_hs__nand3_2 _4311_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1913_),
    .B(_1918_),
    .C(_1922_),
    .Y(_1923_));
 sky130_as_sc_hs__ao22_2 _4312_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1875_),
    .C(_1896_),
    .B(_1894_),
    .D(_1923_),
    .Y(_1924_));
 sky130_as_sc_hs__inv_2 _4313_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_0581_),
    .Y(_1925_));
 sky130_as_sc_hs__nor3_2 _4314_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net38),
    .B(net40),
    .C(_1210_),
    .Y(_1926_));
 sky130_as_sc_hs__ao31_2 _4315_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net38),
    .B(_1162_),
    .C(_1925_),
    .D(_1926_),
    .Y(_1927_));
 sky130_as_sc_hs__nand2_4 _4316_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net48),
    .B(_1927_),
    .Y(_1928_));
 sky130_as_sc_hs__mux2_2 _4317_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1928_),
    .B(net132),
    .A(_0999_),
    .Y(_1929_));
 sky130_as_sc_hs__nand2_2 _4318_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1150_),
    .B(net36),
    .Y(_1930_));
 sky130_as_sc_hs__nand2_2 _4319_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net39),
    .B(_0783_),
    .Y(_1931_));
 sky130_as_sc_hs__nand2_4 _4320_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1930_),
    .B(_1931_),
    .Y(_1932_));
 sky130_as_sc_hs__nand2_4 _4321_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1139_),
    .B(_1932_),
    .Y(_1933_));
 sky130_as_sc_hs__mux2_2 _4322_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1933_),
    .B(_1929_),
    .A(_1924_),
    .Y(_1934_));
 sky130_as_sc_hs__nor2_2 _4323_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net138),
    .B(_1146_),
    .Y(_1935_));
 sky130_as_sc_hs__inv_2 _4324_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_0757_),
    .Y(_1936_));
 sky130_as_sc_hs__oai21_2 _4325_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0656_),
    .B(_1936_),
    .C(_1209_),
    .Y(_1937_));
 sky130_as_sc_hs__nand2_4 _4326_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1935_),
    .B(_1937_),
    .Y(_1938_));
 sky130_as_sc_hs__nor2_2 _4327_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net137),
    .B(_1938_),
    .Y(_1939_));
 sky130_as_sc_hs__nand2_2 _4328_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1934_),
    .B(_1939_),
    .Y(_1940_));
 sky130_as_sc_hs__nand2_2 _4329_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net134),
    .B(\last_A[0] ),
    .Y(_1941_));
 sky130_as_sc_hs__mux2_2 _4330_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1938_),
    .B(_1861_),
    .A(_1941_),
    .Y(_1942_));
 sky130_as_sc_hs__aoi21_2 _4331_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1940_),
    .B(_1942_),
    .C(_1158_),
    .Y(_0399_));
 sky130_as_sc_hs__nand2_2 _4332_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net133),
    .B(_1128_),
    .Y(_1943_));
 sky130_as_sc_hs__nand3_2 _4333_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(carry),
    .B(_1902_),
    .C(_1943_),
    .Y(_1944_));
 sky130_as_sc_hs__nand2_2 _4334_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1861_),
    .B(net40),
    .Y(_1945_));
 sky130_as_sc_hs__nand2_2 _4335_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1863_),
    .B(_1945_),
    .Y(_1946_));
 sky130_as_sc_hs__oa21_2 _4336_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net17),
    .B(_1946_),
    .C(net47),
    .Y(_1947_));
 sky130_as_sc_hs__aoi21_2 _4337_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0928_),
    .B(_0997_),
    .C(_0998_),
    .Y(_1948_));
 sky130_as_sc_hs__aoi21_2 _4338_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1945_),
    .B(_1943_),
    .C(_1948_),
    .Y(_1949_));
 sky130_as_sc_hs__aoi211_2 _4339_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1947_),
    .C(_1949_),
    .D(_1150_),
    .Y(_1950_),
    .A(_1944_));
 sky130_as_sc_hs__or2_2 _4340_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net38),
    .B(_1133_),
    .Y(_1951_));
 sky130_as_sc_hs__aoi22_2 _4341_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net38),
    .B(_1883_),
    .C(_1888_),
    .D(_1951_),
    .Y(_1952_));
 sky130_as_sc_hs__nor2_2 _4342_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net38),
    .B(_0583_),
    .Y(_1953_));
 sky130_as_sc_hs__nor2_2 _4343_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1883_),
    .B(_1888_),
    .Y(_1954_));
 sky130_as_sc_hs__oai21_2 _4344_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1950_),
    .B(_1953_),
    .C(_1954_),
    .Y(_1955_));
 sky130_as_sc_hs__oai21_2 _4345_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1950_),
    .B(_1952_),
    .C(_1955_),
    .Y(_1956_));
 sky130_as_sc_hs__mux2_2 _4346_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1928_),
    .B(net131),
    .A(_1084_),
    .Y(_1957_));
 sky130_as_sc_hs__mux2_2 _4347_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1933_),
    .B(_1957_),
    .A(_1956_),
    .Y(_1958_));
 sky130_as_sc_hs__mux2_2 _4348_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0656_),
    .B(_1958_),
    .A(\last_A[1] ),
    .Y(_1959_));
 sky130_as_sc_hs__inv_2 _4349_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_1938_),
    .Y(_1960_));
 sky130_as_sc_hs__mux2_2 _4350_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1960_),
    .B(_1959_),
    .A(net131),
    .Y(_1961_));
 sky130_as_sc_hs__and2_2 _4351_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net157),
    .B(_1961_),
    .Y(_1962_));
 sky130_as_sc_hs__buff_2 _4352_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1962_),
    .Y(_0400_));
 sky130_as_sc_hs__and2_2 _4353_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1930_),
    .B(_1931_),
    .Y(_1963_));
 sky130_as_sc_hs__buff_4 _4354_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1963_),
    .Y(_1964_));
 sky130_as_sc_hs__nor2_2 _4355_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net31),
    .B(_1964_),
    .Y(_1965_));
 sky130_as_sc_hs__or2_2 _4356_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0648_),
    .B(_0649_),
    .Y(_1966_));
 sky130_as_sc_hs__nand3_2 _4357_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1966_),
    .B(_1867_),
    .C(_1954_),
    .Y(_1967_));
 sky130_as_sc_hs__nand2_2 _4358_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0651_),
    .B(_1890_),
    .Y(_1968_));
 sky130_as_sc_hs__ao21_2 _4359_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1967_),
    .B(_1968_),
    .C(_1863_),
    .Y(_1969_));
 sky130_as_sc_hs__maj3_4 _4360_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1083_),
    .A(net130),
    .C(_1862_),
    .Y(_1970_));
 sky130_as_sc_hs__aoi211_2 _4361_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1948_),
    .C(_1901_),
    .D(_0648_),
    .Y(_1971_),
    .A(net133));
 sky130_as_sc_hs__nand4_2 _4362_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net132),
    .B(_1855_),
    .C(_1859_),
    .Y(_1972_),
    .D(_1860_));
 sky130_as_sc_hs__nor2_2 _4363_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net130),
    .B(_0648_),
    .Y(_1973_));
 sky130_as_sc_hs__oa21_2 _4364_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1083_),
    .B(_1972_),
    .C(_1973_),
    .Y(_1974_));
 sky130_as_sc_hs__aoi211_2 _4365_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1970_),
    .C(_1971_),
    .D(_1974_),
    .Y(_1975_),
    .A(_1128_));
 sky130_as_sc_hs__xnor2_2 _4366_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1882_),
    .Y(_1976_),
    .B(_1975_));
 sky130_as_sc_hs__xnor2_2 _4367_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1969_),
    .Y(_1977_),
    .B(_1976_));
 sky130_as_sc_hs__xnor2_2 _4368_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1906_),
    .Y(_1978_),
    .B(_1970_));
 sky130_as_sc_hs__nor2_2 _4369_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1150_),
    .B(net43),
    .Y(_1979_));
 sky130_as_sc_hs__nor2_2 _4370_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1211_),
    .B(_1906_),
    .Y(_1980_));
 sky130_as_sc_hs__ao21_2 _4371_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1978_),
    .B(_1979_),
    .C(_1980_),
    .Y(_1981_));
 sky130_as_sc_hs__nand2_2 _4372_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1182_),
    .B(_1981_),
    .Y(_1982_));
 sky130_as_sc_hs__nor2_2 _4373_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net37),
    .B(_1123_),
    .Y(_1983_));
 sky130_as_sc_hs__nand2_2 _4374_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net128),
    .B(_1983_),
    .Y(_1984_));
 sky130_as_sc_hs__nand2_2 _4375_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net37),
    .B(_1182_),
    .Y(_1985_));
 sky130_as_sc_hs__xnor2_2 _4376_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1882_),
    .Y(_1986_),
    .B(_1903_));
 sky130_as_sc_hs__oa22_2 _4377_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1094_),
    .B(_1984_),
    .C(_1985_),
    .D(_1986_),
    .Y(_1987_));
 sky130_as_sc_hs__or2_2 _4378_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1129_),
    .B(_1987_),
    .Y(_1988_));
 sky130_as_sc_hs__iao211_2 _4379_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0649_),
    .B(_1977_),
    .C(_1982_),
    .D(_1988_),
    .Y(_1989_));
 sky130_as_sc_hs__inv_2 _4380_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net129),
    .Y(_1990_));
 sky130_as_sc_hs__mux2_2 _4381_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1928_),
    .B(_1990_),
    .A(_1094_),
    .Y(_1991_));
 sky130_as_sc_hs__nor2_2 _4382_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1965_),
    .B(_1991_),
    .Y(_1992_));
 sky130_as_sc_hs__ao21_2 _4383_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1965_),
    .B(_1989_),
    .C(_1992_),
    .Y(_1993_));
 sky130_as_sc_hs__mux2_2 _4384_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1159_),
    .B(_1993_),
    .A(\last_A[2] ),
    .Y(_1994_));
 sky130_as_sc_hs__or2_2 _4385_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1156_),
    .B(_1938_),
    .Y(_1995_));
 sky130_as_sc_hs__inv_2 _4386_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_1995_),
    .Y(_1996_));
 sky130_as_sc_hs__nor2_2 _4387_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1990_),
    .B(_1157_),
    .Y(_1997_));
 sky130_as_sc_hs__ao22_2 _4388_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1994_),
    .C(_1997_),
    .B(_1996_),
    .D(_1938_),
    .Y(_1998_));
 sky130_as_sc_hs__buff_2 _4389_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1998_),
    .Y(_0401_));
 sky130_as_sc_hs__nor2_2 _4390_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1151_),
    .B(_1182_),
    .Y(_1999_));
 sky130_as_sc_hs__aoi21_2 _4391_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1967_),
    .B(_1968_),
    .C(_1863_),
    .Y(_2000_));
 sky130_as_sc_hs__nor2_2 _4392_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net130),
    .B(_0650_),
    .Y(_2001_));
 sky130_as_sc_hs__inv_2 _4393_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_2001_),
    .Y(_2002_));
 sky130_as_sc_hs__nand2_2 _4394_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net130),
    .B(_0651_),
    .Y(_2003_));
 sky130_as_sc_hs__nand3_2 _4395_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1084_),
    .B(_2002_),
    .C(_2003_),
    .Y(_2004_));
 sky130_as_sc_hs__aoi21_2 _4396_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1861_),
    .B(_2002_),
    .C(net17),
    .Y(_2005_));
 sky130_as_sc_hs__oai21_2 _4397_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1861_),
    .B(_0650_),
    .C(\A[1] ),
    .Y(_2006_));
 sky130_as_sc_hs__aoi21_2 _4398_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2002_),
    .B(_2006_),
    .C(_1084_),
    .Y(_2007_));
 sky130_as_sc_hs__aoi21_2 _4399_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2004_),
    .B(_2005_),
    .C(_2007_),
    .Y(_2008_));
 sky130_as_sc_hs__xnor2_2 _4400_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1906_),
    .Y(_2009_),
    .B(_2008_));
 sky130_as_sc_hs__nand2_2 _4401_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2000_),
    .B(_2009_),
    .Y(_2010_));
 sky130_as_sc_hs__nor2_2 _4402_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1990_),
    .B(_1094_),
    .Y(_2011_));
 sky130_as_sc_hs__nor2_2 _4403_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net128),
    .B(_1966_),
    .Y(_2012_));
 sky130_as_sc_hs__maj3_2 _4404_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1084_),
    .A(_1887_),
    .C(_1972_),
    .Y(_2013_));
 sky130_as_sc_hs__oai21_2 _4405_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2011_),
    .B(_2012_),
    .C(_2013_),
    .Y(_2014_));
 sky130_as_sc_hs__or2_2 _4406_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1990_),
    .B(_0650_),
    .Y(_2015_));
 sky130_as_sc_hs__inv_2 _4407_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_2015_),
    .Y(_2016_));
 sky130_as_sc_hs__oai21_2 _4408_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2012_),
    .B(_2016_),
    .C(_0647_),
    .Y(_2017_));
 sky130_as_sc_hs__nor2_2 _4409_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net128),
    .B(_1094_),
    .Y(_2018_));
 sky130_as_sc_hs__oai21_2 _4410_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2018_),
    .B(_2016_),
    .C(_1970_),
    .Y(_2019_));
 sky130_as_sc_hs__nand4_2 _4411_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1910_),
    .B(_2014_),
    .C(_2017_),
    .Y(_2020_),
    .D(_2019_));
 sky130_as_sc_hs__ao31_2 _4412_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2014_),
    .B(_2017_),
    .C(_2019_),
    .D(_1910_),
    .Y(_2021_));
 sky130_as_sc_hs__and2_2 _4413_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2020_),
    .B(_2021_),
    .Y(_2022_));
 sky130_as_sc_hs__xnor2_2 _4414_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2010_),
    .Y(_2023_),
    .B(_2022_));
 sky130_as_sc_hs__maj3_2 _4415_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1094_),
    .A(net128),
    .C(_1903_),
    .Y(_2024_));
 sky130_as_sc_hs__xnor2_2 _4416_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1910_),
    .Y(_2025_),
    .B(_2024_));
 sky130_as_sc_hs__nand2_2 _4417_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\A[3] ),
    .B(_1983_),
    .Y(_2026_));
 sky130_as_sc_hs__oai22_2 _4418_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1985_),
    .B(_2025_),
    .C(_2026_),
    .D(_0754_),
    .Y(_2027_));
 sky130_as_sc_hs__maj3_2 _4419_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_0647_),
    .A(net129),
    .C(_1970_),
    .Y(_2028_));
 sky130_as_sc_hs__xnor2_2 _4420_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1881_),
    .Y(_2029_),
    .B(_2028_));
 sky130_as_sc_hs__nor2_2 _4421_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1211_),
    .B(_1910_),
    .Y(_2030_));
 sky130_as_sc_hs__ao21_2 _4422_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1979_),
    .B(_2029_),
    .C(_2030_),
    .Y(_2031_));
 sky130_as_sc_hs__ao22_2 _4423_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net40),
    .C(_2031_),
    .B(_2027_),
    .D(_1182_),
    .Y(_2032_));
 sky130_as_sc_hs__aoi21_2 _4424_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1999_),
    .B(_2023_),
    .C(_2032_),
    .Y(_2033_));
 sky130_as_sc_hs__mux2_2 _4425_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1928_),
    .B(_1880_),
    .A(_0754_),
    .Y(_2034_));
 sky130_as_sc_hs__mux2_2 _4426_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1933_),
    .B(_2034_),
    .A(_2033_),
    .Y(_2035_));
 sky130_as_sc_hs__nor2_2 _4427_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1159_),
    .B(\last_A[3] ),
    .Y(_2036_));
 sky130_as_sc_hs__mux2_2 _4428_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1938_),
    .B(_1880_),
    .A(_2036_),
    .Y(_2037_));
 sky130_as_sc_hs__buff_8 _4429_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1156_),
    .Y(_2038_));
 sky130_as_sc_hs__aoi211_2 _4430_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2035_),
    .C(_2037_),
    .D(_2038_),
    .Y(_0402_),
    .A(_1939_));
 sky130_as_sc_hs__nand4_2 _4431_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2000_),
    .B(_2009_),
    .C(_2020_),
    .Y(_2039_),
    .D(_2021_));
 sky130_as_sc_hs__or2_2 _4432_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0651_),
    .B(_1879_),
    .Y(_2040_));
 sky130_as_sc_hs__nand2_2 _4433_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1966_),
    .B(_1879_),
    .Y(_2041_));
 sky130_as_sc_hs__nand2_2 _4434_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1880_),
    .B(_0753_),
    .Y(_2042_));
 sky130_as_sc_hs__iao211_2 _4435_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0647_),
    .B(_1970_),
    .C(_2042_),
    .D(net129),
    .Y(_2043_));
 sky130_as_sc_hs__nor2_2 _4436_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1880_),
    .B(_0754_),
    .Y(_2044_));
 sky130_as_sc_hs__aoi31_2 _4437_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0647_),
    .B(_2042_),
    .C(_1970_),
    .D(_2044_),
    .Y(_2045_));
 sky130_as_sc_hs__nand2_2 _4438_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2043_),
    .B(_2045_),
    .Y(_2046_));
 sky130_as_sc_hs__mux2_2 _4439_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2046_),
    .B(_2041_),
    .A(_2040_),
    .Y(_2047_));
 sky130_as_sc_hs__nand2_2 _4440_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0651_),
    .B(_1879_),
    .Y(_2048_));
 sky130_as_sc_hs__or2_2 _4441_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1966_),
    .B(_1879_),
    .Y(_2049_));
 sky130_as_sc_hs__aoi21b_2 _4442_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1900_),
    .B(_1905_),
    .C(_1891_),
    .Y(_2050_));
 sky130_as_sc_hs__mux2_2 _4443_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2050_),
    .B(_2049_),
    .A(_2048_),
    .Y(_2051_));
 sky130_as_sc_hs__nand3_2 _4444_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2039_),
    .B(_2047_),
    .C(_2051_),
    .Y(_2052_));
 sky130_as_sc_hs__ao21_2 _4445_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2047_),
    .B(_2051_),
    .C(_2039_),
    .Y(_2053_));
 sky130_as_sc_hs__nor2_2 _4446_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1151_),
    .B(net46),
    .Y(_2054_));
 sky130_as_sc_hs__nand3_2 _4447_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1128_),
    .B(_2043_),
    .C(_2045_),
    .Y(_2055_));
 sky130_as_sc_hs__ao21_2 _4448_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1899_),
    .B(_1904_),
    .C(_1128_),
    .Y(_2056_));
 sky130_as_sc_hs__inv_2 _4449_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_1879_),
    .Y(_2057_));
 sky130_as_sc_hs__ao21_2 _4450_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2055_),
    .B(_2056_),
    .C(_2057_),
    .Y(_2058_));
 sky130_as_sc_hs__nand3_2 _4451_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2057_),
    .B(_2055_),
    .C(_2056_),
    .Y(_2059_));
 sky130_as_sc_hs__or2_2 _4452_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net46),
    .B(_0840_),
    .Y(_2060_));
 sky130_as_sc_hs__nand2_2 _4453_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net46),
    .B(_1907_),
    .Y(_2061_));
 sky130_as_sc_hs__nand2_2 _4454_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2060_),
    .B(_2061_),
    .Y(_2062_));
 sky130_as_sc_hs__mux2_2 _4455_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net127),
    .B(_2062_),
    .A(_2060_),
    .Y(_2063_));
 sky130_as_sc_hs__nor2_2 _4456_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1211_),
    .B(_2063_),
    .Y(_2064_));
 sky130_as_sc_hs__ao31_2 _4457_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2054_),
    .B(_2058_),
    .C(_2059_),
    .D(_2064_),
    .Y(_2065_));
 sky130_as_sc_hs__aoi31_2 _4458_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1999_),
    .B(_2052_),
    .C(_2053_),
    .D(_2065_),
    .Y(_2066_));
 sky130_as_sc_hs__mux2_2 _4459_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1928_),
    .B(_1244_),
    .A(_1907_),
    .Y(_2067_));
 sky130_as_sc_hs__nor2_2 _4460_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1159_),
    .B(\last_A[4] ),
    .Y(_2068_));
 sky130_as_sc_hs__ao31_2 _4461_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0656_),
    .B(_1933_),
    .C(_2067_),
    .D(_2068_),
    .Y(_2069_));
 sky130_as_sc_hs__aoi21_2 _4462_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1965_),
    .B(_2066_),
    .C(_2069_),
    .Y(_2070_));
 sky130_as_sc_hs__nor2_2 _4463_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1156_),
    .B(_1960_),
    .Y(_2071_));
 sky130_as_sc_hs__ao22_2 _4464_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1996_),
    .C(_2071_),
    .B(_2070_),
    .D(net126),
    .Y(_2072_));
 sky130_as_sc_hs__buff_2 _4465_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2072_),
    .Y(_0403_));
 sky130_as_sc_hs__nand2_2 _4466_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net134),
    .B(\last_A[5] ),
    .Y(_2073_));
 sky130_as_sc_hs__buff_4 _4467_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0918_),
    .Y(_2074_));
 sky130_as_sc_hs__mux2_2 _4468_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1928_),
    .B(net124),
    .A(_2074_),
    .Y(_2075_));
 sky130_as_sc_hs__oai21_2 _4469_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1965_),
    .B(_2075_),
    .C(_1159_),
    .Y(_2076_));
 sky130_as_sc_hs__aoi21_2 _4470_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2073_),
    .B(_2076_),
    .C(_1995_),
    .Y(_2077_));
 sky130_as_sc_hs__clkbuff_4 _4471_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1876_),
    .Y(_2078_));
 sky130_as_sc_hs__nor2_2 _4472_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net127),
    .B(_0651_),
    .Y(_2079_));
 sky130_as_sc_hs__iao211_2 _4473_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1877_),
    .B(_2079_),
    .C(_2045_),
    .D(_2043_),
    .Y(_2080_));
 sky130_as_sc_hs__nand2_2 _4474_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1244_),
    .B(_0840_),
    .Y(_2081_));
 sky130_as_sc_hs__ao31_2 _4475_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1881_),
    .B(_1882_),
    .C(_1889_),
    .D(_2081_),
    .Y(_2082_));
 sky130_as_sc_hs__nand2_2 _4476_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net127),
    .B(_0651_),
    .Y(_2083_));
 sky130_as_sc_hs__ao31_2 _4477_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1881_),
    .B(_1882_),
    .C(_1890_),
    .D(_2083_),
    .Y(_2084_));
 sky130_as_sc_hs__ao22_2 _4478_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1900_),
    .C(_2082_),
    .B(_1905_),
    .D(_2084_),
    .Y(_2085_));
 sky130_as_sc_hs__ao21b_2 _4479_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2079_),
    .B(_2083_),
    .C(_0841_),
    .Y(_2086_));
 sky130_as_sc_hs__nand3_2 _4480_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2080_),
    .B(_2085_),
    .C(_2086_),
    .Y(_2087_));
 sky130_as_sc_hs__xnor2_2 _4481_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2078_),
    .Y(_2088_),
    .B(_2087_));
 sky130_as_sc_hs__xnor2_2 _4482_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2053_),
    .Y(_2089_),
    .B(_2088_));
 sky130_as_sc_hs__nand3_2 _4483_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net125),
    .B(_2074_),
    .C(_1983_),
    .Y(_2090_));
 sky130_as_sc_hs__or2_2 _4484_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1878_),
    .B(_1985_),
    .Y(_2091_));
 sky130_as_sc_hs__or2_2 _4485_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1905_),
    .B(_2091_),
    .Y(_2092_));
 sky130_as_sc_hs__or2_2 _4486_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2078_),
    .B(_2092_),
    .Y(_2093_));
 sky130_as_sc_hs__ao21_2 _4487_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2090_),
    .B(_2093_),
    .C(_1129_),
    .Y(_2094_));
 sky130_as_sc_hs__ao21_2 _4488_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2043_),
    .B(_2045_),
    .C(_1907_),
    .Y(_2095_));
 sky130_as_sc_hs__ao31_2 _4489_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0840_),
    .B(_2043_),
    .C(_2045_),
    .D(_1244_),
    .Y(_2096_));
 sky130_as_sc_hs__nand3_2 _4490_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2078_),
    .B(_2095_),
    .C(_2096_),
    .Y(_2097_));
 sky130_as_sc_hs__ao21_2 _4491_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2095_),
    .B(_2096_),
    .C(_2078_),
    .Y(_2098_));
 sky130_as_sc_hs__nor2_2 _4492_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1211_),
    .B(_2078_),
    .Y(_2099_));
 sky130_as_sc_hs__ao31_2 _4493_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1979_),
    .B(_2097_),
    .C(_2098_),
    .D(_2099_),
    .Y(_2100_));
 sky130_as_sc_hs__ao21_2 _4494_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1900_),
    .B(_1905_),
    .C(_0842_),
    .Y(_2101_));
 sky130_as_sc_hs__ao31_2 _4495_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0842_),
    .B(_1900_),
    .C(_1905_),
    .D(_1244_),
    .Y(_2102_));
 sky130_as_sc_hs__nand3_2 _4496_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2078_),
    .B(_2101_),
    .C(_2102_),
    .Y(_2103_));
 sky130_as_sc_hs__maj3_2 _4497_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_0842_),
    .A(_1244_),
    .C(_1900_),
    .Y(_2104_));
 sky130_as_sc_hs__or2_2 _4498_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2078_),
    .B(_2104_),
    .Y(_2105_));
 sky130_as_sc_hs__aoi211_2 _4499_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2105_),
    .C(_1151_),
    .D(_1129_),
    .Y(_2106_),
    .A(_2103_));
 sky130_as_sc_hs__oai21_2 _4500_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2100_),
    .B(_2106_),
    .C(_1182_),
    .Y(_2107_));
 sky130_as_sc_hs__iao211_2 _4501_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0649_),
    .B(_2089_),
    .C(_2094_),
    .D(_2107_),
    .Y(_2108_));
 sky130_as_sc_hs__ao22_2 _4502_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net124),
    .C(_2077_),
    .B(_2071_),
    .D(_1933_),
    .Y(_2109_));
 sky130_as_sc_hs__ao21_2 _4503_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2077_),
    .B(_2108_),
    .C(_2109_),
    .Y(_2110_));
 sky130_as_sc_hs__buff_2 _4504_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2110_),
    .Y(_0404_));
 sky130_as_sc_hs__mux2_2 _4505_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0757_),
    .B(\last_B[0] ),
    .A(net131),
    .Y(_2111_));
 sky130_as_sc_hs__and2_2 _4506_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net134),
    .B(_2111_),
    .Y(_2112_));
 sky130_as_sc_hs__ao31_2 _4507_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(compat),
    .B(_1139_),
    .C(_1133_),
    .D(_0658_),
    .Y(_2113_));
 sky130_as_sc_hs__and2_2 _4508_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0584_),
    .B(_2113_),
    .Y(_2114_));
 sky130_as_sc_hs__nor2_2 _4509_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net28),
    .B(_1168_),
    .Y(_2115_));
 sky130_as_sc_hs__ao21_2 _4510_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net44),
    .B(_2115_),
    .C(_0660_),
    .Y(_2116_));
 sky130_as_sc_hs__nand2_2 _4511_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net136),
    .B(_2116_),
    .Y(_2117_));
 sky130_as_sc_hs__aoi21_2 _4512_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1209_),
    .B(_2117_),
    .C(_0664_),
    .Y(_2118_));
 sky130_as_sc_hs__oa21_2 _4513_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1209_),
    .B(_2114_),
    .C(_2118_),
    .Y(_2119_));
 sky130_as_sc_hs__buff_4 _4514_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2119_),
    .Y(_2120_));
 sky130_as_sc_hs__mux2_2 _4515_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2120_),
    .B(_2112_),
    .A(\B[0] ),
    .Y(_2121_));
 sky130_as_sc_hs__nor2_2 _4516_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1924_),
    .B(_1964_),
    .Y(_2122_));
 sky130_as_sc_hs__and2_2 _4517_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1159_),
    .B(_2119_),
    .Y(_2123_));
 sky130_as_sc_hs__nand2_2 _4518_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1861_),
    .B(_1964_),
    .Y(_2124_));
 sky130_as_sc_hs__nand2_2 _4519_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2123_),
    .B(_2124_),
    .Y(_2125_));
 sky130_as_sc_hs__nor2_2 _4520_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2122_),
    .B(_2125_),
    .Y(_2126_));
 sky130_as_sc_hs__oa21_2 _4521_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2121_),
    .B(_2126_),
    .C(net149),
    .Y(_2127_));
 sky130_as_sc_hs__buff_2 _4522_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2127_),
    .Y(_0405_));
 sky130_as_sc_hs__mux2_2 _4523_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1932_),
    .B(_1956_),
    .A(net130),
    .Y(_2128_));
 sky130_as_sc_hs__mux2_2 _4524_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_0757_),
    .B(\last_B[1] ),
    .A(net129),
    .Y(_2129_));
 sky130_as_sc_hs__mux2_2 _4525_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net134),
    .B(_2129_),
    .A(_2128_),
    .Y(_2130_));
 sky130_as_sc_hs__mux2_2 _4526_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2120_),
    .B(_2130_),
    .A(\B[1] ),
    .Y(_2131_));
 sky130_as_sc_hs__and2_2 _4527_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net149),
    .B(_2131_),
    .Y(_2132_));
 sky130_as_sc_hs__buff_2 _4528_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2132_),
    .Y(_0406_));
 sky130_as_sc_hs__aoi21_2 _4529_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1990_),
    .B(_1964_),
    .C(net134),
    .Y(_2133_));
 sky130_as_sc_hs__oai21_2 _4530_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1964_),
    .B(_1989_),
    .C(_2133_),
    .Y(_2134_));
 sky130_as_sc_hs__buff_8 _4531_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0757_),
    .Y(_2135_));
 sky130_as_sc_hs__mux2_2 _4532_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2135_),
    .B(\last_B[2] ),
    .A(\A[3] ),
    .Y(_2136_));
 sky130_as_sc_hs__nand2_2 _4533_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net134),
    .B(_2136_),
    .Y(_2137_));
 sky130_as_sc_hs__oai21_2 _4534_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net166),
    .B(_2120_),
    .C(net150),
    .Y(_2138_));
 sky130_as_sc_hs__aoi31_2 _4535_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2120_),
    .B(_2134_),
    .C(_2137_),
    .D(net167),
    .Y(_0407_));
 sky130_as_sc_hs__ao21_2 _4536_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1880_),
    .B(_1964_),
    .C(net137),
    .Y(_2139_));
 sky130_as_sc_hs__ao21_2 _4537_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1932_),
    .B(_2033_),
    .C(_2139_),
    .Y(_2140_));
 sky130_as_sc_hs__mux2_2 _4538_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2135_),
    .B(\last_B[3] ),
    .A(net126),
    .Y(_2141_));
 sky130_as_sc_hs__nand2_2 _4539_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net134),
    .B(_2141_),
    .Y(_2142_));
 sky130_as_sc_hs__oai21_2 _4540_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net169),
    .B(_2120_),
    .C(net150),
    .Y(_2143_));
 sky130_as_sc_hs__aoi31_2 _4541_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2120_),
    .B(_2140_),
    .C(_2142_),
    .D(_2143_),
    .Y(_0408_));
 sky130_as_sc_hs__mux2_2 _4542_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1932_),
    .B(_2066_),
    .A(_1244_),
    .Y(_2144_));
 sky130_as_sc_hs__mux2_2 _4543_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2135_),
    .B(\last_B[4] ),
    .A(net124),
    .Y(_2145_));
 sky130_as_sc_hs__nor2_2 _4544_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1159_),
    .B(_2145_),
    .Y(_2146_));
 sky130_as_sc_hs__mux2_2 _4545_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2120_),
    .B(_2146_),
    .A(_1243_),
    .Y(_2147_));
 sky130_as_sc_hs__aoi211_2 _4546_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2144_),
    .C(_2147_),
    .D(_2038_),
    .Y(_0409_),
    .A(_2123_));
 sky130_as_sc_hs__nand2_2 _4547_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1932_),
    .B(_2123_),
    .Y(_2148_));
 sky130_as_sc_hs__ao21_2 _4548_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_B[5] ),
    .B(_0757_),
    .C(_0656_),
    .Y(_2149_));
 sky130_as_sc_hs__ao31_2 _4549_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(carry),
    .B(_1133_),
    .C(_2115_),
    .D(_2149_),
    .Y(_2150_));
 sky130_as_sc_hs__mux2_2 _4550_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2119_),
    .B(_2150_),
    .A(\B[5] ),
    .Y(_2151_));
 sky130_as_sc_hs__nand2_2 _4551_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net157),
    .B(_2151_),
    .Y(_2152_));
 sky130_as_sc_hs__aoi31_2 _4552_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1919_),
    .B(_1964_),
    .C(_2123_),
    .D(_2152_),
    .Y(_2153_));
 sky130_as_sc_hs__oa21_2 _4553_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2108_),
    .B(_2148_),
    .C(_2153_),
    .Y(_2154_));
 sky130_as_sc_hs__buff_2 _4554_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2154_),
    .Y(_0410_));
 sky130_as_sc_hs__nand2_2 _4555_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2095_),
    .B(_2096_),
    .Y(_2155_));
 sky130_as_sc_hs__maj3_2 _4556_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2074_),
    .A(net125),
    .C(_2155_),
    .Y(_2156_));
 sky130_as_sc_hs__nor2_2 _4557_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net43),
    .B(_2156_),
    .Y(_2157_));
 sky130_as_sc_hs__nor2_2 _4558_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1129_),
    .B(_1923_),
    .Y(_2158_));
 sky130_as_sc_hs__oai22_2 _4559_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2053_),
    .B(_2088_),
    .C(_2157_),
    .D(_2158_),
    .Y(_2159_));
 sky130_as_sc_hs__oai21_2 _4560_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1001_),
    .B(_1930_),
    .C(_1931_),
    .Y(_2160_));
 sky130_as_sc_hs__nand2_2 _4561_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0656_),
    .B(_2160_),
    .Y(_2161_));
 sky130_as_sc_hs__oai21_2 _4562_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1169_),
    .B(_1002_),
    .C(net133),
    .Y(_2162_));
 sky130_as_sc_hs__nor2_2 _4563_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0577_),
    .B(_1895_),
    .Y(_2163_));
 sky130_as_sc_hs__aoi21_2 _4564_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1169_),
    .B(_2163_),
    .C(net133),
    .Y(_2164_));
 sky130_as_sc_hs__aoi21_2 _4565_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1139_),
    .B(_2162_),
    .C(_2164_),
    .Y(_2165_));
 sky130_as_sc_hs__mux2_2 _4566_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1936_),
    .B(_2165_),
    .A(\last_flags[0] ),
    .Y(_2166_));
 sky130_as_sc_hs__nand3_2 _4567_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net135),
    .B(_1925_),
    .C(_2163_),
    .Y(_2167_));
 sky130_as_sc_hs__ao31_2 _4568_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\instr_cycle[1] ),
    .B(_0783_),
    .C(_2113_),
    .D(net135),
    .Y(_2168_));
 sky130_as_sc_hs__nand4_2 _4569_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1935_),
    .B(_1127_),
    .C(_2167_),
    .Y(_2169_),
    .D(_2168_));
 sky130_as_sc_hs__aoi21_2 _4570_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net135),
    .B(_2166_),
    .C(_2169_),
    .Y(_2170_));
 sky130_as_sc_hs__ao21_2 _4571_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1863_),
    .B(_2169_),
    .C(_1130_),
    .Y(_2171_));
 sky130_as_sc_hs__ao21_2 _4572_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2161_),
    .B(_2170_),
    .C(_2171_),
    .Y(_2172_));
 sky130_as_sc_hs__nor2_2 _4573_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0649_),
    .B(_2172_),
    .Y(_2173_));
 sky130_as_sc_hs__ao31_2 _4574_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2074_),
    .B(_2101_),
    .C(_2102_),
    .D(_1919_),
    .Y(_2174_));
 sky130_as_sc_hs__ao21_2 _4575_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2101_),
    .B(_2102_),
    .C(_2074_),
    .Y(_2175_));
 sky130_as_sc_hs__nand3_2 _4576_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net43),
    .B(_2174_),
    .C(_2175_),
    .Y(_2176_));
 sky130_as_sc_hs__iao211_2 _4577_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net43),
    .B(_2156_),
    .C(_2176_),
    .D(_2054_),
    .Y(_2177_));
 sky130_as_sc_hs__aoi21_2 _4578_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2170_),
    .B(_2177_),
    .C(_2172_),
    .Y(_2178_));
 sky130_as_sc_hs__ao21_2 _4579_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2159_),
    .B(_2173_),
    .C(_2178_),
    .Y(_2179_));
 sky130_as_sc_hs__buff_2 _4580_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2179_),
    .Y(_0411_));
 sky130_as_sc_hs__nor2_2 _4581_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net126),
    .B(\A[3] ),
    .Y(_2180_));
 sky130_as_sc_hs__nand4_2 _4582_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1919_),
    .B(_1990_),
    .C(_1887_),
    .Y(_2181_),
    .D(_2180_));
 sky130_as_sc_hs__ao31_2 _4583_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(carry),
    .B(_1133_),
    .C(_2115_),
    .D(_2181_),
    .Y(_2182_));
 sky130_as_sc_hs__nand2_2 _4584_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\last_flags[1] ),
    .B(_2135_),
    .Y(_2183_));
 sky130_as_sc_hs__iao211_2 _4585_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2135_),
    .B(_2182_),
    .C(_2183_),
    .D(net135),
    .Y(_2184_));
 sky130_as_sc_hs__mux2_2 _4586_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2118_),
    .B(_2184_),
    .A(zero),
    .Y(_2185_));
 sky130_as_sc_hs__nand2_2 _4587_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net160),
    .B(_2185_),
    .Y(_2186_));
 sky130_as_sc_hs__nand2_2 _4588_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0652_),
    .B(_1896_),
    .Y(_2187_));
 sky130_as_sc_hs__or2_2 _4589_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(compat),
    .B(_2187_),
    .Y(_2188_));
 sky130_as_sc_hs__nor3_2 _4590_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0647_),
    .B(_0999_),
    .C(_2188_),
    .Y(_2189_));
 sky130_as_sc_hs__nand4_2 _4591_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0754_),
    .B(_1907_),
    .C(_1901_),
    .Y(_2190_),
    .D(_2189_));
 sky130_as_sc_hs__ao31_2 _4592_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net42),
    .B(_0652_),
    .C(_1983_),
    .D(zero),
    .Y(_2191_));
 sky130_as_sc_hs__aoi22_2 _4593_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(compat),
    .B(_2191_),
    .C(_2187_),
    .D(zero),
    .Y(_2192_));
 sky130_as_sc_hs__oai21_2 _4594_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2074_),
    .B(_2190_),
    .C(_2192_),
    .Y(_2193_));
 sky130_as_sc_hs__oai21_2 _4595_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2124_),
    .B(_2181_),
    .C(_2114_),
    .Y(_2194_));
 sky130_as_sc_hs__aoi21b_2 _4596_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\instr_cycle[1] ),
    .B(_1935_),
    .C(zero),
    .Y(_2195_));
 sky130_as_sc_hs__aoi211_2 _4597_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2194_),
    .C(net135),
    .D(_2195_),
    .Y(_2196_),
    .A(_2193_));
 sky130_as_sc_hs__nor3_2 _4598_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1956_),
    .B(_1989_),
    .C(_2186_),
    .Y(_2197_));
 sky130_as_sc_hs__nand4_2 _4599_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2033_),
    .B(_2066_),
    .C(_2122_),
    .Y(_2198_),
    .D(_2197_));
 sky130_as_sc_hs__oai22_2 _4600_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2186_),
    .B(_2196_),
    .C(_2198_),
    .D(_2108_),
    .Y(_0412_));
 sky130_as_sc_hs__inv_2 _4601_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[0] ),
    .Y(_2199_));
 sky130_as_sc_hs__clkbuff_4 _4602_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0534_),
    .Y(_2200_));
 sky130_as_sc_hs__inv_2 _4603_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(in_irupt),
    .Y(_2201_));
 sky130_as_sc_hs__nand3_2 _4604_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2201_),
    .B(net138),
    .C(needs_irupt),
    .Y(_2202_));
 sky130_as_sc_hs__oa21_2 _4605_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net138),
    .B(_1143_),
    .C(_2202_),
    .Y(_2203_));
 sky130_as_sc_hs__and2_2 _4606_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0657_),
    .B(_0660_),
    .Y(_2204_));
 sky130_as_sc_hs__buff_2 _4607_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2204_),
    .Y(_2205_));
 sky130_as_sc_hs__ao22_2 _4608_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2199_),
    .C(_2205_),
    .B(_2203_),
    .D(\last_PC[0] ),
    .Y(_2206_));
 sky130_as_sc_hs__aoi21_2 _4609_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2200_),
    .B(_0999_),
    .C(_2206_),
    .Y(_2207_));
 sky130_as_sc_hs__iao211_2 _4610_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1150_),
    .B(_1162_),
    .C(_1286_),
    .D(_1930_),
    .Y(_2208_));
 sky130_as_sc_hs__mux2_2 _4611_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_1138_),
    .B(_1001_),
    .A(net42),
    .Y(_2209_));
 sky130_as_sc_hs__ao22_2 _4612_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net30),
    .C(_2209_),
    .B(_2208_),
    .D(_1000_),
    .Y(_2210_));
 sky130_as_sc_hs__aoi31_2 _4613_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(zero),
    .B(_1123_),
    .C(net41),
    .D(net32),
    .Y(_2211_));
 sky130_as_sc_hs__ao31_2 _4614_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(carry),
    .B(net32),
    .C(net41),
    .D(_2211_),
    .Y(_2212_));
 sky130_as_sc_hs__oai21_2 _4615_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(zero),
    .B(net44),
    .C(_1139_),
    .Y(_2213_));
 sky130_as_sc_hs__aoi211_2 _4616_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2213_),
    .C(_1209_),
    .D(_0584_),
    .Y(_2214_),
    .A(net47));
 sky130_as_sc_hs__nand2_2 _4617_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net32),
    .B(_2163_),
    .Y(_2215_));
 sky130_as_sc_hs__aoi22_2 _4618_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2212_),
    .B(_2214_),
    .C(_2215_),
    .D(net136),
    .Y(_2216_));
 sky130_as_sc_hs__aoi21_2 _4619_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1143_),
    .B(_2210_),
    .C(_2216_),
    .Y(_2217_));
 sky130_as_sc_hs__oa21_2 _4620_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net139),
    .B(_2217_),
    .C(_0533_),
    .Y(_2218_));
 sky130_as_sc_hs__clkbuff_4 _4621_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2218_),
    .Y(_2219_));
 sky130_as_sc_hs__mux2_2 _4622_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2219_),
    .B(_2207_),
    .A(_2199_),
    .Y(_2220_));
 sky130_as_sc_hs__nor2_2 _4623_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1180_),
    .B(_2220_),
    .Y(_0413_));
 sky130_as_sc_hs__inv_2 _4624_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[1] ),
    .Y(_2221_));
 sky130_as_sc_hs__xnor2_2 _4625_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2221_),
    .Y(_2222_),
    .B(\PC[0] ));
 sky130_as_sc_hs__buff_2 _4626_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2203_),
    .Y(_2223_));
 sky130_as_sc_hs__ao22_2 _4627_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_PC[1] ),
    .C(_2222_),
    .B(_2205_),
    .D(_2223_),
    .Y(_2224_));
 sky130_as_sc_hs__aoi21_2 _4628_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2200_),
    .B(_1084_),
    .C(_2224_),
    .Y(_2225_));
 sky130_as_sc_hs__buff_2 _4629_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2218_),
    .Y(_2226_));
 sky130_as_sc_hs__mux2_2 _4630_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2226_),
    .B(_2225_),
    .A(_2221_),
    .Y(_2227_));
 sky130_as_sc_hs__nor2_2 _4631_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1180_),
    .B(_2227_),
    .Y(_0414_));
 sky130_as_sc_hs__nor2_2 _4632_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2221_),
    .B(_2199_),
    .Y(_2228_));
 sky130_as_sc_hs__xnor2_2 _4633_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[2] ),
    .Y(_2229_),
    .B(_2228_));
 sky130_as_sc_hs__nor2_2 _4634_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2135_),
    .B(_2229_),
    .Y(_2230_));
 sky130_as_sc_hs__ao31_2 _4635_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0663_),
    .B(\last_PC[2] ),
    .C(_2135_),
    .D(_2230_),
    .Y(_2231_));
 sky130_as_sc_hs__clkbuff_4 _4636_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2202_),
    .Y(_2232_));
 sky130_as_sc_hs__oai21_2 _4637_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0663_),
    .B(_2229_),
    .C(_2232_),
    .Y(_2233_));
 sky130_as_sc_hs__ao21_2 _4638_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net135),
    .B(_2231_),
    .C(_2233_),
    .Y(_2234_));
 sky130_as_sc_hs__aoi21_2 _4639_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2200_),
    .B(_0647_),
    .C(_2234_),
    .Y(_2235_));
 sky130_as_sc_hs__oai21_2 _4640_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net182),
    .B(_2219_),
    .C(net160),
    .Y(_2236_));
 sky130_as_sc_hs__aoi21_2 _4641_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2219_),
    .B(_2235_),
    .C(_2236_),
    .Y(_0415_));
 sky130_as_sc_hs__inv_2 _4642_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[3] ),
    .Y(_2237_));
 sky130_as_sc_hs__or2_2 _4643_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net139),
    .B(net135),
    .Y(_2238_));
 sky130_as_sc_hs__nand2_2 _4644_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\PC[2] ),
    .B(_2228_),
    .Y(_2239_));
 sky130_as_sc_hs__xnor2_2 _4645_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[3] ),
    .Y(_2240_),
    .B(_2239_));
 sky130_as_sc_hs__aoi22_2 _4646_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_PC[3] ),
    .B(_2205_),
    .C(_2240_),
    .D(_2223_),
    .Y(_2241_));
 sky130_as_sc_hs__oa21_2 _4647_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2238_),
    .B(_0754_),
    .C(_2241_),
    .Y(_2242_));
 sky130_as_sc_hs__mux2_2 _4648_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2226_),
    .B(_2242_),
    .A(_2237_),
    .Y(_2243_));
 sky130_as_sc_hs__nor2_2 _4649_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1180_),
    .B(_2243_),
    .Y(_0416_));
 sky130_as_sc_hs__inv_2 _4650_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[4] ),
    .Y(_2244_));
 sky130_as_sc_hs__nor2_2 _4651_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2237_),
    .B(_2239_),
    .Y(_2245_));
 sky130_as_sc_hs__xnor2_2 _4652_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2244_),
    .Y(_2246_),
    .B(_2245_));
 sky130_as_sc_hs__ao22_2 _4653_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_PC[4] ),
    .C(_2246_),
    .B(_2205_),
    .D(_2223_),
    .Y(_2247_));
 sky130_as_sc_hs__aoi21_2 _4654_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2200_),
    .B(_0842_),
    .C(_2247_),
    .Y(_2248_));
 sky130_as_sc_hs__nor2_2 _4655_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\PC[4] ),
    .B(_2219_),
    .Y(_2249_));
 sky130_as_sc_hs__aoi211_2 _4656_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2248_),
    .C(_2249_),
    .D(_2038_),
    .Y(_0417_),
    .A(_2219_));
 sky130_as_sc_hs__nand2_2 _4657_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\PC[4] ),
    .B(_2245_),
    .Y(_2250_));
 sky130_as_sc_hs__xnor2_2 _4658_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[5] ),
    .Y(_2251_),
    .B(_2250_));
 sky130_as_sc_hs__ao22_2 _4659_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\last_PC[5] ),
    .C(_2251_),
    .B(_2205_),
    .D(_2223_),
    .Y(_2252_));
 sky130_as_sc_hs__aoi21_2 _4660_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2200_),
    .B(_2074_),
    .C(_2252_),
    .Y(_2253_));
 sky130_as_sc_hs__nor2_2 _4661_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net592),
    .B(_2219_),
    .Y(_2254_));
 sky130_as_sc_hs__aoi211_2 _4662_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2253_),
    .C(_2254_),
    .D(_2038_),
    .Y(_0418_),
    .A(_2219_));
 sky130_as_sc_hs__buff_2 _4663_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2202_),
    .Y(_2255_));
 sky130_as_sc_hs__oai21_2 _4664_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net138),
    .B(_1143_),
    .C(_2255_),
    .Y(_2256_));
 sky130_as_sc_hs__clkbuff_4 _4665_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2256_),
    .Y(_2257_));
 sky130_as_sc_hs__nand3_2 _4666_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\PC[5] ),
    .B(\PC[4] ),
    .C(_2245_),
    .Y(_2258_));
 sky130_as_sc_hs__inv_2 _4667_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_2258_),
    .Y(_2259_));
 sky130_as_sc_hs__clkbuff_4 _4668_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2218_),
    .Y(_2260_));
 sky130_as_sc_hs__oai21_2 _4669_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2257_),
    .B(_2259_),
    .C(_2260_),
    .Y(_2261_));
 sky130_as_sc_hs__inv_2 _4670_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[6] ),
    .Y(_2262_));
 sky130_as_sc_hs__ao22_2 _4671_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[0] ),
    .C(_2205_),
    .B(_2200_),
    .D(\last_PC[6] ),
    .Y(_2263_));
 sky130_as_sc_hs__ao31_2 _4672_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2262_),
    .B(_2223_),
    .C(_2259_),
    .D(_2263_),
    .Y(_2264_));
 sky130_as_sc_hs__ao22_2 _4673_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[6] ),
    .C(_2264_),
    .B(_2261_),
    .D(_2226_),
    .Y(_2265_));
 sky130_as_sc_hs__and2_2 _4674_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net158),
    .B(_2265_),
    .Y(_2266_));
 sky130_as_sc_hs__buff_2 _4675_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2266_),
    .Y(_0419_));
 sky130_as_sc_hs__nor2_2 _4676_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2262_),
    .B(_2258_),
    .Y(_2267_));
 sky130_as_sc_hs__oai21_2 _4677_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2257_),
    .B(_2267_),
    .C(_2260_),
    .Y(_2268_));
 sky130_as_sc_hs__inv_2 _4678_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[7] ),
    .Y(_2269_));
 sky130_as_sc_hs__ao22_2 _4679_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[1] ),
    .C(_2205_),
    .B(_2200_),
    .D(\last_PC[7] ),
    .Y(_2270_));
 sky130_as_sc_hs__ao31_2 _4680_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2269_),
    .B(_2223_),
    .C(_2267_),
    .D(_2270_),
    .Y(_2271_));
 sky130_as_sc_hs__ao22_2 _4681_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[7] ),
    .C(_2271_),
    .B(_2268_),
    .D(_2226_),
    .Y(_2272_));
 sky130_as_sc_hs__and2_2 _4682_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net158),
    .B(_2272_),
    .Y(_2273_));
 sky130_as_sc_hs__buff_2 _4683_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2273_),
    .Y(_0420_));
 sky130_as_sc_hs__and2_2 _4684_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[7] ),
    .B(_2267_),
    .Y(_2274_));
 sky130_as_sc_hs__oai21_2 _4685_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2257_),
    .B(_2274_),
    .C(_2260_),
    .Y(_2275_));
 sky130_as_sc_hs__inv_2 _4686_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[8] ),
    .Y(_2276_));
 sky130_as_sc_hs__ao22_2 _4687_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[2] ),
    .C(_2204_),
    .B(_0675_),
    .D(\last_PC[8] ),
    .Y(_2277_));
 sky130_as_sc_hs__ao31_2 _4688_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2276_),
    .B(_2203_),
    .C(_2274_),
    .D(_2277_),
    .Y(_2278_));
 sky130_as_sc_hs__ao22_2 _4689_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[8] ),
    .C(_2278_),
    .B(_2275_),
    .D(_2226_),
    .Y(_2279_));
 sky130_as_sc_hs__and2_2 _4690_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net155),
    .B(_2279_),
    .Y(_2280_));
 sky130_as_sc_hs__buff_2 _4691_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2280_),
    .Y(_0421_));
 sky130_as_sc_hs__and2_2 _4692_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[8] ),
    .B(_2274_),
    .Y(_2281_));
 sky130_as_sc_hs__oai21_2 _4693_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2257_),
    .B(_2281_),
    .C(_2260_),
    .Y(_2282_));
 sky130_as_sc_hs__inv_2 _4694_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[9] ),
    .Y(_2283_));
 sky130_as_sc_hs__ao22_2 _4695_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[3] ),
    .C(_2204_),
    .B(_0675_),
    .D(\last_PC[9] ),
    .Y(_2284_));
 sky130_as_sc_hs__ao31_2 _4696_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2283_),
    .B(_2203_),
    .C(_2281_),
    .D(_2284_),
    .Y(_2285_));
 sky130_as_sc_hs__ao22_2 _4697_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[9] ),
    .C(_2285_),
    .B(_2282_),
    .D(_2226_),
    .Y(_2286_));
 sky130_as_sc_hs__and2_2 _4698_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net155),
    .B(_2286_),
    .Y(_2287_));
 sky130_as_sc_hs__buff_2 _4699_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2287_),
    .Y(_0422_));
 sky130_as_sc_hs__and2_2 _4700_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[9] ),
    .B(_2281_),
    .Y(_2288_));
 sky130_as_sc_hs__oai21_2 _4701_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2257_),
    .B(_2288_),
    .C(_2260_),
    .Y(_2289_));
 sky130_as_sc_hs__inv_2 _4702_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[10] ),
    .Y(_2290_));
 sky130_as_sc_hs__ao22_2 _4703_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[4] ),
    .C(_2204_),
    .B(_0675_),
    .D(\last_PC[10] ),
    .Y(_2291_));
 sky130_as_sc_hs__ao31_2 _4704_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2290_),
    .B(_2203_),
    .C(_2288_),
    .D(_2291_),
    .Y(_2292_));
 sky130_as_sc_hs__ao22_2 _4705_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[10] ),
    .C(_2292_),
    .B(_2289_),
    .D(_2226_),
    .Y(_2293_));
 sky130_as_sc_hs__and2_2 _4706_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net155),
    .B(_2293_),
    .Y(_2294_));
 sky130_as_sc_hs__buff_2 _4707_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2294_),
    .Y(_0423_));
 sky130_as_sc_hs__ao21_2 _4708_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[10] ),
    .B(_2288_),
    .C(_2256_),
    .Y(_2295_));
 sky130_as_sc_hs__nand2_2 _4709_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2260_),
    .B(_2295_),
    .Y(_2296_));
 sky130_as_sc_hs__nor2_2 _4710_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\PC[11] ),
    .B(_2290_),
    .Y(_2297_));
 sky130_as_sc_hs__ao22_2 _4711_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\P[5] ),
    .C(_2204_),
    .B(_0675_),
    .D(\last_PC[11] ),
    .Y(_2298_));
 sky130_as_sc_hs__ao31_2 _4712_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2223_),
    .B(_2288_),
    .C(_2297_),
    .D(_2298_),
    .Y(_2299_));
 sky130_as_sc_hs__ao22_2 _4713_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[11] ),
    .C(_2299_),
    .B(_2296_),
    .D(_2260_),
    .Y(_2300_));
 sky130_as_sc_hs__and2_2 _4714_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net158),
    .B(_2300_),
    .Y(_2301_));
 sky130_as_sc_hs__buff_2 _4715_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2301_),
    .Y(_0424_));
 sky130_as_sc_hs__nor2_2 _4716_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0665_),
    .B(_2167_),
    .Y(_2302_));
 sky130_as_sc_hs__xnor2_2 _4717_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net584),
    .Y(_2303_),
    .B(_2302_));
 sky130_as_sc_hs__nand2_2 _4718_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net160),
    .B(_2303_),
    .Y(_0425_));
 sky130_as_sc_hs__nand4_2 _4719_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net150),
    .B(\ROM_dest[1] ),
    .C(_0532_),
    .Y(_2304_),
    .D(_1011_));
 sky130_as_sc_hs__mux2_2 _4720_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2304_),
    .B(net256),
    .A(\ROM_spi_dat_out[0] ),
    .Y(_2305_));
 sky130_as_sc_hs__buff_2 _4721_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2305_),
    .Y(_0426_));
 sky130_as_sc_hs__mux2_2 _4722_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2304_),
    .B(net184),
    .A(\ROM_spi_dat_out[1] ),
    .Y(_2306_));
 sky130_as_sc_hs__buff_2 _4723_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2306_),
    .Y(_0427_));
 sky130_as_sc_hs__mux2_2 _4724_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2304_),
    .B(net175),
    .A(\ROM_spi_dat_out[2] ),
    .Y(_2307_));
 sky130_as_sc_hs__buff_2 _4725_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2307_),
    .Y(_0428_));
 sky130_as_sc_hs__mux2_2 _4726_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2304_),
    .B(net589),
    .A(\ROM_spi_dat_out[3] ),
    .Y(_2308_));
 sky130_as_sc_hs__buff_2 _4727_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2308_),
    .Y(_0429_));
 sky130_as_sc_hs__mux2_2 _4728_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2304_),
    .B(net591),
    .A(\ROM_spi_dat_out[4] ),
    .Y(_2309_));
 sky130_as_sc_hs__buff_2 _4729_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2309_),
    .Y(_0430_));
 sky130_as_sc_hs__mux2_2 _4730_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2304_),
    .B(net579),
    .A(\ROM_spi_dat_out[5] ),
    .Y(_2310_));
 sky130_as_sc_hs__buff_2 _4731_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2310_),
    .Y(_0431_));
 sky130_as_sc_hs__nor2_2 _4732_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1146_),
    .B(_2202_),
    .Y(_2311_));
 sky130_as_sc_hs__and2_2 _4733_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net154),
    .B(_2311_),
    .Y(_2312_));
 sky130_as_sc_hs__buff_4 _4734_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2312_),
    .Y(_2313_));
 sky130_as_sc_hs__buff_4 _4735_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2313_),
    .Y(_2314_));
 sky130_as_sc_hs__mux2_2 _4736_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2314_),
    .B(\PC[0] ),
    .A(net406),
    .Y(_2315_));
 sky130_as_sc_hs__buff_2 _4737_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net407),
    .Y(_0432_));
 sky130_as_sc_hs__mux2_2 _4738_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2314_),
    .B(\PC[1] ),
    .A(net460),
    .Y(_2316_));
 sky130_as_sc_hs__buff_2 _4739_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net461),
    .Y(_0433_));
 sky130_as_sc_hs__mux2_2 _4740_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2314_),
    .B(\PC[2] ),
    .A(net205),
    .Y(_2317_));
 sky130_as_sc_hs__buff_2 _4741_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2317_),
    .Y(_0434_));
 sky130_as_sc_hs__mux2_2 _4742_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2314_),
    .B(\PC[3] ),
    .A(net574),
    .Y(_2318_));
 sky130_as_sc_hs__buff_2 _4743_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net575),
    .Y(_0435_));
 sky130_as_sc_hs__mux2_2 _4744_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2314_),
    .B(\PC[4] ),
    .A(net417),
    .Y(_2319_));
 sky130_as_sc_hs__buff_2 _4745_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2319_),
    .Y(_0436_));
 sky130_as_sc_hs__mux2_2 _4746_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2314_),
    .B(\PC[5] ),
    .A(net221),
    .Y(_2320_));
 sky130_as_sc_hs__buff_2 _4747_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2320_),
    .Y(_0437_));
 sky130_as_sc_hs__mux2_2 _4748_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2314_),
    .B(\PC[6] ),
    .A(net186),
    .Y(_2321_));
 sky130_as_sc_hs__buff_2 _4749_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net187),
    .Y(_0438_));
 sky130_as_sc_hs__buff_8 _4750_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2313_),
    .Y(_2322_));
 sky130_as_sc_hs__mux2_2 _4751_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2322_),
    .B(\PC[7] ),
    .A(net185),
    .Y(_2323_));
 sky130_as_sc_hs__buff_2 _4752_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2323_),
    .Y(_0439_));
 sky130_as_sc_hs__mux2_2 _4753_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2322_),
    .B(\PC[8] ),
    .A(net183),
    .Y(_2324_));
 sky130_as_sc_hs__buff_2 _4754_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2324_),
    .Y(_0440_));
 sky130_as_sc_hs__mux2_2 _4755_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2322_),
    .B(\PC[9] ),
    .A(net181),
    .Y(_2325_));
 sky130_as_sc_hs__buff_2 _4756_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2325_),
    .Y(_0441_));
 sky130_as_sc_hs__mux2_2 _4757_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2322_),
    .B(\PC[10] ),
    .A(net176),
    .Y(_2326_));
 sky130_as_sc_hs__buff_2 _4758_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2326_),
    .Y(_0442_));
 sky130_as_sc_hs__mux2_2 _4759_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2322_),
    .B(\PC[11] ),
    .A(net178),
    .Y(_2327_));
 sky130_as_sc_hs__buff_2 _4760_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2327_),
    .Y(_0443_));
 sky130_as_sc_hs__mux2_2 _4761_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2322_),
    .B(carry),
    .A(net564),
    .Y(_2328_));
 sky130_as_sc_hs__buff_2 _4762_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2328_),
    .Y(_0444_));
 sky130_as_sc_hs__mux2_2 _4763_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2322_),
    .B(zero),
    .A(net556),
    .Y(_2329_));
 sky130_as_sc_hs__buff_2 _4764_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2329_),
    .Y(_0445_));
 sky130_as_sc_hs__buff_4 _4765_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2313_),
    .Y(_2330_));
 sky130_as_sc_hs__mux2_2 _4766_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2330_),
    .B(net132),
    .A(net560),
    .Y(_2331_));
 sky130_as_sc_hs__buff_2 _4767_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2331_),
    .Y(_0446_));
 sky130_as_sc_hs__mux2_2 _4768_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2330_),
    .B(net131),
    .A(net220),
    .Y(_2332_));
 sky130_as_sc_hs__buff_2 _4769_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2332_),
    .Y(_0447_));
 sky130_as_sc_hs__mux2_2 _4770_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2330_),
    .B(net129),
    .A(net286),
    .Y(_2333_));
 sky130_as_sc_hs__buff_2 _4771_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2333_),
    .Y(_0448_));
 sky130_as_sc_hs__mux2_2 _4772_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2330_),
    .B(\A[3] ),
    .A(net566),
    .Y(_2334_));
 sky130_as_sc_hs__buff_2 _4773_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2334_),
    .Y(_0449_));
 sky130_as_sc_hs__mux2_2 _4774_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2330_),
    .B(net126),
    .A(net582),
    .Y(_2335_));
 sky130_as_sc_hs__buff_2 _4775_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2335_),
    .Y(_0450_));
 sky130_as_sc_hs__mux2_2 _4776_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2330_),
    .B(net124),
    .A(net570),
    .Y(_2336_));
 sky130_as_sc_hs__buff_2 _4777_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2336_),
    .Y(_0451_));
 sky130_as_sc_hs__mux2_2 _4778_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2330_),
    .B(\B[0] ),
    .A(net533),
    .Y(_2337_));
 sky130_as_sc_hs__buff_2 _4779_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net534),
    .Y(_0452_));
 sky130_as_sc_hs__buff_4 _4780_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2313_),
    .Y(_2338_));
 sky130_as_sc_hs__mux2_2 _4781_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2338_),
    .B(\B[1] ),
    .A(net500),
    .Y(_2339_));
 sky130_as_sc_hs__buff_2 _4782_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net501),
    .Y(_0453_));
 sky130_as_sc_hs__mux2_2 _4783_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2338_),
    .B(net166),
    .A(net206),
    .Y(_2340_));
 sky130_as_sc_hs__buff_2 _4784_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2340_),
    .Y(_0454_));
 sky130_as_sc_hs__mux2_2 _4785_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2338_),
    .B(net169),
    .A(net219),
    .Y(_2341_));
 sky130_as_sc_hs__buff_2 _4786_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2341_),
    .Y(_0455_));
 sky130_as_sc_hs__mux2_2 _4787_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2338_),
    .B(\B[4] ),
    .A(net448),
    .Y(_2342_));
 sky130_as_sc_hs__buff_2 _4788_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net449),
    .Y(_0456_));
 sky130_as_sc_hs__mux2_2 _4789_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2338_),
    .B(\B[5] ),
    .A(net212),
    .Y(_2343_));
 sky130_as_sc_hs__buff_2 _4790_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net213),
    .Y(_0457_));
 sky130_as_sc_hs__mux2_2 _4791_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2338_),
    .B(net122),
    .A(net443),
    .Y(_2344_));
 sky130_as_sc_hs__buff_2 _4792_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2344_),
    .Y(_0458_));
 sky130_as_sc_hs__mux2_2 _4793_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2338_),
    .B(net102),
    .A(net367),
    .Y(_2345_));
 sky130_as_sc_hs__buff_2 _4794_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2345_),
    .Y(_0459_));
 sky130_as_sc_hs__buff_4 _4795_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2312_),
    .Y(_2346_));
 sky130_as_sc_hs__mux2_2 _4796_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2346_),
    .B(net61),
    .A(net189),
    .Y(_2347_));
 sky130_as_sc_hs__buff_2 _4797_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2347_),
    .Y(_0460_));
 sky130_as_sc_hs__mux2_2 _4798_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2346_),
    .B(net53),
    .A(net174),
    .Y(_2348_));
 sky130_as_sc_hs__buff_2 _4799_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2348_),
    .Y(_0461_));
 sky130_as_sc_hs__mux2_2 _4800_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2346_),
    .B(net50),
    .A(net333),
    .Y(_2349_));
 sky130_as_sc_hs__buff_2 _4801_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2349_),
    .Y(_0462_));
 sky130_as_sc_hs__mux2_2 _4802_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2346_),
    .B(net142),
    .A(net245),
    .Y(_2350_));
 sky130_as_sc_hs__buff_2 _4803_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2350_),
    .Y(_0463_));
 sky130_as_sc_hs__mux2_2 _4804_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2346_),
    .B(\P[0] ),
    .A(net180),
    .Y(_2351_));
 sky130_as_sc_hs__buff_2 _4805_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2351_),
    .Y(_0464_));
 sky130_as_sc_hs__mux2_2 _4806_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2346_),
    .B(\P[1] ),
    .A(net392),
    .Y(_2352_));
 sky130_as_sc_hs__buff_2 _4807_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2352_),
    .Y(_0465_));
 sky130_as_sc_hs__mux2_2 _4808_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2346_),
    .B(\P[2] ),
    .A(net190),
    .Y(_2353_));
 sky130_as_sc_hs__buff_2 _4809_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2353_),
    .Y(_0466_));
 sky130_as_sc_hs__mux2_2 _4810_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2313_),
    .B(\P[3] ),
    .A(net177),
    .Y(_2354_));
 sky130_as_sc_hs__buff_2 _4811_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2354_),
    .Y(_0467_));
 sky130_as_sc_hs__mux2_2 _4812_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2313_),
    .B(\P[4] ),
    .A(net201),
    .Y(_2355_));
 sky130_as_sc_hs__buff_2 _4813_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2355_),
    .Y(_0468_));
 sky130_as_sc_hs__mux2_2 _4814_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2313_),
    .B(\P[5] ),
    .A(net194),
    .Y(_2356_));
 sky130_as_sc_hs__buff_2 _4815_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2356_),
    .Y(_0469_));
 sky130_as_sc_hs__inv_2 _4816_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(last_inter),
    .Y(_2357_));
 sky130_as_sc_hs__aoi21_2 _4817_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net16),
    .B(_2357_),
    .C(net172),
    .Y(_2358_));
 sky130_as_sc_hs__nor3_2 _4818_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1157_),
    .B(_2311_),
    .C(net173),
    .Y(_0470_));
 sky130_as_sc_hs__ao31_2 _4819_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net136),
    .B(_0761_),
    .C(_2257_),
    .D(_2201_),
    .Y(_2359_));
 sky130_as_sc_hs__nand3_2 _4820_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net138),
    .B(_0761_),
    .C(_2257_),
    .Y(_2360_));
 sky130_as_sc_hs__aoi21_2 _4821_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2359_),
    .B(_2360_),
    .C(_1158_),
    .Y(_0471_));
 sky130_as_sc_hs__nand3_2 _4822_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net143),
    .B(\mem_cycle[1] ),
    .C(net144),
    .Y(_2361_));
 sky130_as_sc_hs__oai21_2 _4823_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(spi_clkdiv),
    .B(net8),
    .C(_0530_),
    .Y(_2362_));
 sky130_as_sc_hs__inv_2 _4824_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_2362_),
    .Y(_2363_));
 sky130_as_sc_hs__ao31_4 _4825_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0668_),
    .B(_0531_),
    .C(_2361_),
    .D(_2363_),
    .Y(_2364_));
 sky130_as_sc_hs__or2_2 _4826_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[0] ),
    .B(_2364_),
    .Y(_2365_));
 sky130_as_sc_hs__nand2_4 _4827_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[0] ),
    .B(_2364_),
    .Y(_2366_));
 sky130_as_sc_hs__nand3_2 _4828_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net146),
    .B(_2365_),
    .C(_2366_),
    .Y(_2367_));
 sky130_as_sc_hs__inv_2 _4829_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_2367_),
    .Y(_0472_));
 sky130_as_sc_hs__or2_2 _4830_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[1] ),
    .B(_2366_),
    .Y(_2368_));
 sky130_as_sc_hs__ao21_2 _4831_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[4] ),
    .B(_0527_),
    .C(_2368_),
    .Y(_2369_));
 sky130_as_sc_hs__nand2_2 _4832_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net586),
    .B(_2366_),
    .Y(_2370_));
 sky130_as_sc_hs__aoi21_2 _4833_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2369_),
    .B(_2370_),
    .C(_1158_),
    .Y(_0473_));
 sky130_as_sc_hs__nor2_2 _4834_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_0526_),
    .B(_2366_),
    .Y(_2371_));
 sky130_as_sc_hs__xnor2_2 _4835_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net577),
    .Y(_2372_),
    .B(_2371_));
 sky130_as_sc_hs__nor2_2 _4836_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1180_),
    .B(_2372_),
    .Y(_0474_));
 sky130_as_sc_hs__nand2_2 _4837_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\ROM_spi_cycle[2] ),
    .B(\ROM_spi_cycle[1] ),
    .Y(_2373_));
 sky130_as_sc_hs__nand2_2 _4838_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\ROM_spi_cycle[3] ),
    .B(\ROM_spi_cycle[0] ),
    .Y(_2374_));
 sky130_as_sc_hs__and2_2 _4839_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[4] ),
    .B(\ROM_spi_cycle[0] ),
    .Y(_2375_));
 sky130_as_sc_hs__oai21_2 _4840_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0529_),
    .B(_2375_),
    .C(_0528_),
    .Y(_2376_));
 sky130_as_sc_hs__oai21_2 _4841_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2373_),
    .B(_2374_),
    .C(_2376_),
    .Y(_2377_));
 sky130_as_sc_hs__nor2_2 _4842_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2366_),
    .B(_2373_),
    .Y(_2378_));
 sky130_as_sc_hs__nor2_2 _4843_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\ROM_spi_cycle[3] ),
    .B(_2378_),
    .Y(_2379_));
 sky130_as_sc_hs__aoi211_2 _4844_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2377_),
    .C(_2379_),
    .D(_1735_),
    .Y(_0475_),
    .A(_2364_));
 sky130_as_sc_hs__or2_2 _4845_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[2] ),
    .B(_2368_),
    .Y(_2380_));
 sky130_as_sc_hs__ao21_2 _4846_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[4] ),
    .B(_2380_),
    .C(\ROM_spi_cycle[3] ),
    .Y(_2381_));
 sky130_as_sc_hs__aoi31_2 _4847_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[4] ),
    .B(\ROM_spi_cycle[3] ),
    .C(_2378_),
    .D(_2038_),
    .Y(_2382_));
 sky130_as_sc_hs__iao211_2 _4848_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net571),
    .B(_2378_),
    .C(_2381_),
    .D(_2382_),
    .Y(_2383_));
 sky130_as_sc_hs__inv_2 _4849_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(_2383_),
    .Y(_0476_));
 sky130_as_sc_hs__and2_2 _4850_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net152),
    .B(net16),
    .Y(_2384_));
 sky130_as_sc_hs__buff_2 _4851_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2384_),
    .Y(_0477_));
 sky130_as_sc_hs__nor2_2 _4852_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net143),
    .B(_1292_),
    .Y(_2385_));
 sky130_as_sc_hs__inv_2 _4853_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(CS_ROM),
    .Y(_2386_));
 sky130_as_sc_hs__ao31_2 _4854_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1284_),
    .B(_1354_),
    .C(_2385_),
    .D(_2386_),
    .Y(_2387_));
 sky130_as_sc_hs__nand2_2 _4855_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\mem_cycle[1] ),
    .B(_2387_),
    .Y(_2388_));
 sky130_as_sc_hs__ao31_2 _4856_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net144),
    .B(_1354_),
    .C(_2385_),
    .D(CS_ROM),
    .Y(_2389_));
 sky130_as_sc_hs__ao21_2 _4857_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2388_),
    .B(_2389_),
    .C(_1735_),
    .Y(_2390_));
 sky130_as_sc_hs__buff_2 _4858_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2390_),
    .Y(_0478_));
 sky130_as_sc_hs__or2_2 _4859_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[0] ),
    .B(_2362_),
    .Y(_2391_));
 sky130_as_sc_hs__nor2_4 _4860_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1297_),
    .B(_0531_),
    .Y(_2392_));
 sky130_as_sc_hs__buff_8 _4861_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2392_),
    .Y(_2393_));
 sky130_as_sc_hs__nand2_2 _4862_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(SCLK_ROM),
    .B(_2362_),
    .Y(_2394_));
 sky130_as_sc_hs__ao21_2 _4863_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1354_),
    .B(_2393_),
    .C(_2394_),
    .Y(_2395_));
 sky130_as_sc_hs__aoi21_2 _4864_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2391_),
    .B(_2395_),
    .C(_1158_),
    .Y(_0479_));
 sky130_as_sc_hs__mux2_2 _4865_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2366_),
    .B(ROM_DO),
    .A(\ROM_spi_dat_out[7] ),
    .Y(_2396_));
 sky130_as_sc_hs__and2_2 _4866_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net148),
    .B(_2396_),
    .Y(_2397_));
 sky130_as_sc_hs__buff_2 _4867_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2397_),
    .Y(_0480_));
 sky130_as_sc_hs__oai21_2 _4868_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_cycle[0] ),
    .B(_2362_),
    .C(_2364_),
    .Y(_2398_));
 sky130_as_sc_hs__clkbuff_4 _4869_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2398_),
    .Y(_2399_));
 sky130_as_sc_hs__nand2_2 _4870_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1296_),
    .B(net144),
    .Y(_2400_));
 sky130_as_sc_hs__oai22_2 _4871_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_addr_buff[8] ),
    .B(net145),
    .C(_2400_),
    .D(\ROM_addr_buff[0] ),
    .Y(_2401_));
 sky130_as_sc_hs__xnor2_2 _4872_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net143),
    .Y(_2402_),
    .B(net144));
 sky130_as_sc_hs__nor2_2 _4873_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_1296_),
    .B(_2402_),
    .Y(_2403_));
 sky130_as_sc_hs__aoi211_2 _4874_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2401_),
    .C(_2403_),
    .D(_1293_),
    .Y(_2404_),
    .A(\mem_cycle[2] ));
 sky130_as_sc_hs__aoi211_2 _4875_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1293_),
    .C(_2399_),
    .D(_2404_),
    .Y(_2405_),
    .A(net9));
 sky130_as_sc_hs__aoi211_2 _4876_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2399_),
    .C(_2405_),
    .D(_1735_),
    .Y(_0481_),
    .A(_1181_));
 sky130_as_sc_hs__oai22_2 _4877_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net27),
    .B(net145),
    .C(_2400_),
    .D(\ROM_addr_buff[1] ),
    .Y(_2406_));
 sky130_as_sc_hs__aoi211_2 _4878_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2406_),
    .C(_2403_),
    .D(_1293_),
    .Y(_2407_),
    .A(\mem_cycle[2] ));
 sky130_as_sc_hs__aoi211_2 _4879_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_1293_),
    .C(_2399_),
    .D(_2407_),
    .Y(_2408_),
    .A(\ROM_spi_dat_out[0] ));
 sky130_as_sc_hs__aoi211_2 _4880_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .B(_2399_),
    .C(_2408_),
    .D(_1735_),
    .Y(_0482_),
    .A(_1187_));
 sky130_as_sc_hs__inv_2 _4881_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(net143),
    .Y(_2409_));
 sky130_as_sc_hs__nor2_2 _4882_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2409_),
    .B(\mem_cycle[1] ),
    .Y(_2410_));
 sky130_as_sc_hs__mux2_2 _4883_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net145),
    .B(\ROM_addr_buff[2] ),
    .A(\ROM_addr_buff[10] ),
    .Y(_2411_));
 sky130_as_sc_hs__and2_2 _4884_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_dat_out[1] ),
    .B(_1292_),
    .Y(_2412_));
 sky130_as_sc_hs__ao31_2 _4885_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1285_),
    .B(_2410_),
    .C(_2411_),
    .D(_2412_),
    .Y(_2413_));
 sky130_as_sc_hs__mux2_2 _4886_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2399_),
    .B(\ROM_spi_dat_out[2] ),
    .A(_2413_),
    .Y(_2414_));
 sky130_as_sc_hs__and2_2 _4887_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net151),
    .B(_2414_),
    .Y(_2415_));
 sky130_as_sc_hs__buff_2 _4888_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2415_),
    .Y(_0483_));
 sky130_as_sc_hs__mux2_2 _4889_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(net145),
    .B(\ROM_addr_buff[3] ),
    .A(\ROM_addr_buff[11] ),
    .Y(_2416_));
 sky130_as_sc_hs__and2_2 _4890_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_dat_out[2] ),
    .B(_1292_),
    .Y(_2417_));
 sky130_as_sc_hs__ao31_2 _4891_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1285_),
    .B(_2410_),
    .C(_2416_),
    .D(_2417_),
    .Y(_2418_));
 sky130_as_sc_hs__mux2_2 _4892_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2399_),
    .B(\ROM_spi_dat_out[3] ),
    .A(_2418_),
    .Y(_2419_));
 sky130_as_sc_hs__and2_2 _4893_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net151),
    .B(_2419_),
    .Y(_2420_));
 sky130_as_sc_hs__buff_2 _4894_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2420_),
    .Y(_0484_));
 sky130_as_sc_hs__nor2_2 _4895_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2409_),
    .B(_2400_),
    .Y(_2421_));
 sky130_as_sc_hs__and2_2 _4896_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_dat_out[3] ),
    .B(_1292_),
    .Y(_2422_));
 sky130_as_sc_hs__ao31_2 _4897_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_addr_buff[4] ),
    .B(_1285_),
    .C(_2421_),
    .D(_2422_),
    .Y(_2423_));
 sky130_as_sc_hs__mux2_2 _4898_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2399_),
    .B(\ROM_spi_dat_out[4] ),
    .A(_2423_),
    .Y(_2424_));
 sky130_as_sc_hs__and2_2 _4899_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net151),
    .B(_2424_),
    .Y(_2425_));
 sky130_as_sc_hs__buff_2 _4900_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2425_),
    .Y(_0485_));
 sky130_as_sc_hs__and2_2 _4901_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_dat_out[4] ),
    .B(_1292_),
    .Y(_2426_));
 sky130_as_sc_hs__ao31_2 _4902_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_addr_buff[5] ),
    .B(_1285_),
    .C(_2421_),
    .D(_2426_),
    .Y(_2427_));
 sky130_as_sc_hs__mux2_2 _4903_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2398_),
    .B(\ROM_spi_dat_out[5] ),
    .A(_2427_),
    .Y(_2428_));
 sky130_as_sc_hs__and2_2 _4904_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net151),
    .B(_2428_),
    .Y(_2429_));
 sky130_as_sc_hs__buff_2 _4905_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2429_),
    .Y(_0486_));
 sky130_as_sc_hs__and2_2 _4906_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_dat_out[5] ),
    .B(_1292_),
    .Y(_2430_));
 sky130_as_sc_hs__ao31_2 _4907_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_addr_buff[6] ),
    .B(_1285_),
    .C(_2421_),
    .D(_2430_),
    .Y(_2431_));
 sky130_as_sc_hs__mux2_2 _4908_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2398_),
    .B(\ROM_spi_dat_out[6] ),
    .A(_2431_),
    .Y(_2432_));
 sky130_as_sc_hs__and2_2 _4909_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net151),
    .B(_2432_),
    .Y(_2433_));
 sky130_as_sc_hs__buff_2 _4910_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2433_),
    .Y(_0487_));
 sky130_as_sc_hs__and2_2 _4911_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_spi_dat_out[6] ),
    .B(_0530_),
    .Y(_2434_));
 sky130_as_sc_hs__ao31_2 _4912_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\ROM_addr_buff[7] ),
    .B(_1285_),
    .C(_2421_),
    .D(_2434_),
    .Y(_2435_));
 sky130_as_sc_hs__mux2_2 _4913_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2398_),
    .B(\ROM_spi_dat_out[7] ),
    .A(_2435_),
    .Y(_2436_));
 sky130_as_sc_hs__and2_2 _4914_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net152),
    .B(_2436_),
    .Y(_2437_));
 sky130_as_sc_hs__buff_2 _4915_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2437_),
    .Y(_0488_));
 sky130_as_sc_hs__and2_2 _4916_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[0] ),
    .B(_2232_),
    .Y(_2438_));
 sky130_as_sc_hs__nand2_4 _4917_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_0533_),
    .B(_1290_),
    .Y(_2439_));
 sky130_as_sc_hs__buff_4 _4918_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2439_),
    .Y(_2440_));
 sky130_as_sc_hs__mux2_2 _4919_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2440_),
    .B(\ROM_addr_buff[0] ),
    .A(_2438_),
    .Y(_2441_));
 sky130_as_sc_hs__and2_2 _4920_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net159),
    .B(_2441_),
    .Y(_2442_));
 sky130_as_sc_hs__buff_2 _4921_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2442_),
    .Y(_0489_));
 sky130_as_sc_hs__and2_2 _4922_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[1] ),
    .B(_2232_),
    .Y(_2443_));
 sky130_as_sc_hs__mux2_2 _4923_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2440_),
    .B(\ROM_addr_buff[1] ),
    .A(_2443_),
    .Y(_2444_));
 sky130_as_sc_hs__and2_2 _4924_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net159),
    .B(_2444_),
    .Y(_2445_));
 sky130_as_sc_hs__buff_2 _4925_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2445_),
    .Y(_0490_));
 sky130_as_sc_hs__nand2_2 _4926_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(net593),
    .B(_2440_),
    .Y(_2446_));
 sky130_as_sc_hs__inv_2 _4927_ (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(\PC[2] ),
    .Y(_2447_));
 sky130_as_sc_hs__ao21_2 _4928_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2447_),
    .B(_2232_),
    .C(_2440_),
    .Y(_2448_));
 sky130_as_sc_hs__aoi21_2 _4929_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_2446_),
    .B(_2448_),
    .C(_1158_),
    .Y(_0491_));
 sky130_as_sc_hs__and2_2 _4930_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[3] ),
    .B(_2232_),
    .Y(_2449_));
 sky130_as_sc_hs__mux2_2 _4931_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2440_),
    .B(\ROM_addr_buff[3] ),
    .A(_2449_),
    .Y(_2450_));
 sky130_as_sc_hs__and2_2 _4932_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net159),
    .B(_2450_),
    .Y(_2451_));
 sky130_as_sc_hs__buff_2 _4933_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2451_),
    .Y(_0492_));
 sky130_as_sc_hs__and2_2 _4934_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[4] ),
    .B(_2232_),
    .Y(_2452_));
 sky130_as_sc_hs__mux2_2 _4935_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2440_),
    .B(\ROM_addr_buff[4] ),
    .A(_2452_),
    .Y(_2453_));
 sky130_as_sc_hs__and2_2 _4936_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net158),
    .B(_2453_),
    .Y(_2454_));
 sky130_as_sc_hs__buff_2 _4937_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2454_),
    .Y(_0493_));
 sky130_as_sc_hs__and2_2 _4938_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[5] ),
    .B(_2255_),
    .Y(_2455_));
 sky130_as_sc_hs__mux2_2 _4939_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2439_),
    .B(\ROM_addr_buff[5] ),
    .A(_2455_),
    .Y(_2456_));
 sky130_as_sc_hs__and2_2 _4940_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net158),
    .B(_2456_),
    .Y(_2457_));
 sky130_as_sc_hs__buff_2 _4941_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2457_),
    .Y(_0494_));
 sky130_as_sc_hs__and2_2 _4942_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[6] ),
    .B(_2255_),
    .Y(_2458_));
 sky130_as_sc_hs__mux2_2 _4943_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2439_),
    .B(\ROM_addr_buff[6] ),
    .A(_2458_),
    .Y(_2459_));
 sky130_as_sc_hs__and2_2 _4944_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net154),
    .B(_2459_),
    .Y(_2460_));
 sky130_as_sc_hs__buff_2 _4945_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2460_),
    .Y(_0495_));
 sky130_as_sc_hs__and2_2 _4946_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[7] ),
    .B(_2255_),
    .Y(_2461_));
 sky130_as_sc_hs__mux2_2 _4947_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2439_),
    .B(\ROM_addr_buff[7] ),
    .A(_2461_),
    .Y(_2462_));
 sky130_as_sc_hs__and2_2 _4948_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net154),
    .B(_2462_),
    .Y(_2463_));
 sky130_as_sc_hs__buff_2 _4949_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2463_),
    .Y(_0496_));
 sky130_as_sc_hs__and2_2 _4950_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[8] ),
    .B(_2255_),
    .Y(_2464_));
 sky130_as_sc_hs__mux2_2 _4951_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2439_),
    .B(\ROM_addr_buff[8] ),
    .A(_2464_),
    .Y(_2465_));
 sky130_as_sc_hs__and2_2 _4952_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net154),
    .B(_2465_),
    .Y(_2466_));
 sky130_as_sc_hs__buff_2 _4953_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2466_),
    .Y(_0497_));
 sky130_as_sc_hs__and2_2 _4954_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[9] ),
    .B(_2255_),
    .Y(_2467_));
 sky130_as_sc_hs__mux2_2 _4955_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2439_),
    .B(net27),
    .A(_2467_),
    .Y(_2468_));
 sky130_as_sc_hs__and2_2 _4956_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net154),
    .B(_2468_),
    .Y(_2469_));
 sky130_as_sc_hs__buff_2 _4957_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2469_),
    .Y(_0498_));
 sky130_as_sc_hs__and2_2 _4958_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(\PC[10] ),
    .B(_2255_),
    .Y(_2470_));
 sky130_as_sc_hs__mux2_2 _4959_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2439_),
    .B(\ROM_addr_buff[10] ),
    .A(_2470_),
    .Y(_2471_));
 sky130_as_sc_hs__and2_2 _4960_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net155),
    .B(_2471_),
    .Y(_2472_));
 sky130_as_sc_hs__buff_2 _4961_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2472_),
    .Y(_0499_));
 sky130_as_sc_hs__nand2_2 _4962_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(\PC[11] ),
    .B(_2232_),
    .Y(_2473_));
 sky130_as_sc_hs__mux2_2 _4963_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2440_),
    .B(_1306_),
    .A(_2473_),
    .Y(_2474_));
 sky130_as_sc_hs__nor2_2 _4964_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2038_),
    .B(_2474_),
    .Y(_0500_));
 sky130_as_sc_hs__mux2_2 _4965_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2393_),
    .B(\ROM_addr_buff[0] ),
    .A(\last_addr[0] ),
    .Y(_2475_));
 sky130_as_sc_hs__and2_2 _4966_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net159),
    .B(_2475_),
    .Y(_2476_));
 sky130_as_sc_hs__buff_2 _4967_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2476_),
    .Y(_0501_));
 sky130_as_sc_hs__mux2_2 _4968_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2393_),
    .B(\ROM_addr_buff[1] ),
    .A(\last_addr[1] ),
    .Y(_2477_));
 sky130_as_sc_hs__and2_2 _4969_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net159),
    .B(_2477_),
    .Y(_2478_));
 sky130_as_sc_hs__buff_2 _4970_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2478_),
    .Y(_0502_));
 sky130_as_sc_hs__mux2_2 _4971_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2393_),
    .B(\ROM_addr_buff[2] ),
    .A(\last_addr[2] ),
    .Y(_2479_));
 sky130_as_sc_hs__and2_2 _4972_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net159),
    .B(_2479_),
    .Y(_2480_));
 sky130_as_sc_hs__buff_2 _4973_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2480_),
    .Y(_0503_));
 sky130_as_sc_hs__mux2_2 _4974_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2393_),
    .B(\ROM_addr_buff[3] ),
    .A(\last_addr[3] ),
    .Y(_2481_));
 sky130_as_sc_hs__and2_2 _4975_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net159),
    .B(_2481_),
    .Y(_2482_));
 sky130_as_sc_hs__buff_2 _4976_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2482_),
    .Y(_0504_));
 sky130_as_sc_hs__mux2_2 _4977_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2393_),
    .B(\ROM_addr_buff[4] ),
    .A(\last_addr[4] ),
    .Y(_2483_));
 sky130_as_sc_hs__and2_2 _4978_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net158),
    .B(_2483_),
    .Y(_2484_));
 sky130_as_sc_hs__buff_2 _4979_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2484_),
    .Y(_0505_));
 sky130_as_sc_hs__mux2_2 _4980_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2393_),
    .B(\ROM_addr_buff[5] ),
    .A(\last_addr[5] ),
    .Y(_2485_));
 sky130_as_sc_hs__and2_2 _4981_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net158),
    .B(_2485_),
    .Y(_2486_));
 sky130_as_sc_hs__buff_2 _4982_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2486_),
    .Y(_0506_));
 sky130_as_sc_hs__mux2_2 _4983_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2392_),
    .B(\ROM_addr_buff[6] ),
    .A(\last_addr[6] ),
    .Y(_2487_));
 sky130_as_sc_hs__and2_2 _4984_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net152),
    .B(_2487_),
    .Y(_2488_));
 sky130_as_sc_hs__buff_2 _4985_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2488_),
    .Y(_0507_));
 sky130_as_sc_hs__mux2_2 _4986_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2392_),
    .B(\ROM_addr_buff[7] ),
    .A(\last_addr[7] ),
    .Y(_2489_));
 sky130_as_sc_hs__and2_2 _4987_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net153),
    .B(_2489_),
    .Y(_2490_));
 sky130_as_sc_hs__buff_2 _4988_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2490_),
    .Y(_0508_));
 sky130_as_sc_hs__mux2_2 _4989_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2392_),
    .B(\ROM_addr_buff[8] ),
    .A(\last_addr[8] ),
    .Y(_2491_));
 sky130_as_sc_hs__and2_2 _4990_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net156),
    .B(_2491_),
    .Y(_2492_));
 sky130_as_sc_hs__buff_2 _4991_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2492_),
    .Y(_0509_));
 sky130_as_sc_hs__mux2_2 _4992_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2392_),
    .B(net27),
    .A(\last_addr[9] ),
    .Y(_2493_));
 sky130_as_sc_hs__and2_2 _4993_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net156),
    .B(_2493_),
    .Y(_2494_));
 sky130_as_sc_hs__buff_2 _4994_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2494_),
    .Y(_0510_));
 sky130_as_sc_hs__mux2_2 _4995_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2392_),
    .B(\ROM_addr_buff[10] ),
    .A(\last_addr[10] ),
    .Y(_2495_));
 sky130_as_sc_hs__and2_2 _4996_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net155),
    .B(_2495_),
    .Y(_2496_));
 sky130_as_sc_hs__buff_2 _4997_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2496_),
    .Y(_0511_));
 sky130_as_sc_hs__mux2_2 _4998_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2392_),
    .B(\ROM_addr_buff[11] ),
    .A(\last_addr[11] ),
    .Y(_2497_));
 sky130_as_sc_hs__and2_2 _4999_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net156),
    .B(_2497_),
    .Y(_2498_));
 sky130_as_sc_hs__buff_2 _5000_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2498_),
    .Y(_0512_));
 sky130_as_sc_hs__xnor2_2 _5001_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(net170),
    .Y(_2499_),
    .B(_1293_));
 sky130_as_sc_hs__nor2_2 _5002_ (.VNB(VGND),
    .VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .A(_2038_),
    .B(net171),
    .Y(_0513_));
 sky130_as_sc_hs__nor2_4 _5003_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1224_),
    .B(_1366_),
    .Y(_2500_));
 sky130_as_sc_hs__mux2_2 _5004_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2500_),
    .B(_1470_),
    .A(net179),
    .Y(_2501_));
 sky130_as_sc_hs__buff_2 _5005_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2501_),
    .Y(_0514_));
 sky130_as_sc_hs__mux2_2 _5006_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2500_),
    .B(_1475_),
    .A(net191),
    .Y(_2502_));
 sky130_as_sc_hs__buff_2 _5007_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2502_),
    .Y(_0515_));
 sky130_as_sc_hs__mux2_2 _5008_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2500_),
    .B(_1478_),
    .A(net193),
    .Y(_2503_));
 sky130_as_sc_hs__buff_2 _5009_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2503_),
    .Y(_0516_));
 sky130_as_sc_hs__mux2_2 _5010_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2500_),
    .B(_1481_),
    .A(net423),
    .Y(_2504_));
 sky130_as_sc_hs__buff_2 _5011_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2504_),
    .Y(_0517_));
 sky130_as_sc_hs__mux2_2 _5012_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2500_),
    .B(_1484_),
    .A(net494),
    .Y(_2505_));
 sky130_as_sc_hs__buff_2 _5013_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2505_),
    .Y(_0518_));
 sky130_as_sc_hs__mux2_2 _5014_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2500_),
    .B(_1487_),
    .A(net518),
    .Y(_2506_));
 sky130_as_sc_hs__buff_2 _5015_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2506_),
    .Y(_0519_));
 sky130_as_sc_hs__nor2_4 _5016_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .A(_1274_),
    .B(_1554_),
    .Y(_2507_));
 sky130_as_sc_hs__mux2_2 _5017_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2507_),
    .B(_1470_),
    .A(net374),
    .Y(_2508_));
 sky130_as_sc_hs__buff_2 _5018_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2508_),
    .Y(_0520_));
 sky130_as_sc_hs__mux2_2 _5019_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2507_),
    .B(_1475_),
    .A(net561),
    .Y(_2509_));
 sky130_as_sc_hs__buff_2 _5020_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2509_),
    .Y(_0521_));
 sky130_as_sc_hs__mux2_2 _5021_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2507_),
    .B(_1478_),
    .A(net345),
    .Y(_2510_));
 sky130_as_sc_hs__buff_2 _5022_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2510_),
    .Y(_0522_));
 sky130_as_sc_hs__mux2_2 _5023_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2507_),
    .B(_1481_),
    .A(net509),
    .Y(_2511_));
 sky130_as_sc_hs__buff_2 _5024_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2511_),
    .Y(_0523_));
 sky130_as_sc_hs__mux2_2 _5025_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2507_),
    .B(_1484_),
    .A(net275),
    .Y(_2512_));
 sky130_as_sc_hs__buff_2 _5026_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2512_),
    .Y(_0524_));
 sky130_as_sc_hs__mux2_2 _5027_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .S(_2507_),
    .B(_1487_),
    .A(net434),
    .Y(_2513_));
 sky130_as_sc_hs__buff_2 _5028_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2513_),
    .Y(_0525_));
 sky130_as_sc_hs__dfxtp_2 _5029_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[44][0] ),
    .D(_0024_));
 sky130_as_sc_hs__dfxtp_2 _5030_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[44][1] ),
    .D(_0025_));
 sky130_as_sc_hs__dfxtp_2 _5031_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[44][2] ),
    .D(_0026_));
 sky130_as_sc_hs__dfxtp_2 _5032_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[44][3] ),
    .D(_0027_));
 sky130_as_sc_hs__dfxtp_2 _5033_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[44][4] ),
    .D(_0028_));
 sky130_as_sc_hs__dfxtp_2 _5034_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[44][5] ),
    .D(_0029_));
 sky130_as_sc_hs__dfxtp_2 _5035_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[45][0] ),
    .D(_0030_));
 sky130_as_sc_hs__dfxtp_2 _5036_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[45][1] ),
    .D(_0031_));
 sky130_as_sc_hs__dfxtp_2 _5037_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(\RAM[45][2] ),
    .D(_0032_));
 sky130_as_sc_hs__dfxtp_2 _5038_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[45][3] ),
    .D(_0033_));
 sky130_as_sc_hs__dfxtp_2 _5039_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[45][4] ),
    .D(_0034_));
 sky130_as_sc_hs__dfxtp_2 _5040_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[45][5] ),
    .D(_0035_));
 sky130_as_sc_hs__dfxtp_2 _5041_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[62][0] ),
    .D(_0036_));
 sky130_as_sc_hs__dfxtp_2 _5042_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\RAM[62][1] ),
    .D(_0037_));
 sky130_as_sc_hs__dfxtp_2 _5043_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[62][2] ),
    .D(_0038_));
 sky130_as_sc_hs__dfxtp_2 _5044_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(\RAM[62][3] ),
    .D(_0039_));
 sky130_as_sc_hs__dfxtp_2 _5045_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[62][4] ),
    .D(_0040_));
 sky130_as_sc_hs__dfxtp_2 _5046_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[62][5] ),
    .D(_0041_));
 sky130_as_sc_hs__dfxtp_2 _5047_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[49][0] ),
    .D(_0042_));
 sky130_as_sc_hs__dfxtp_2 _5048_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[49][1] ),
    .D(_0043_));
 sky130_as_sc_hs__dfxtp_2 _5049_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[49][2] ),
    .D(_0044_));
 sky130_as_sc_hs__dfxtp_2 _5050_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[49][3] ),
    .D(_0045_));
 sky130_as_sc_hs__dfxtp_2 _5051_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[49][4] ),
    .D(_0046_));
 sky130_as_sc_hs__dfxtp_2 _5052_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[49][5] ),
    .D(_0047_));
 sky130_as_sc_hs__dfxtp_2 _5053_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\mem_cycle[0] ),
    .D(_0048_));
 sky130_as_sc_hs__dfxtp_4 _5054_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem_cycle[1] ),
    .D(_0049_));
 sky130_as_sc_hs__dfxtp_2 _5055_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\mem_cycle[2] ),
    .D(_0050_));
 sky130_as_sc_hs__dfxtp_2 _5056_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[46][0] ),
    .D(_0051_));
 sky130_as_sc_hs__dfxtp_2 _5057_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[46][1] ),
    .D(_0052_));
 sky130_as_sc_hs__dfxtp_2 _5058_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[46][2] ),
    .D(_0053_));
 sky130_as_sc_hs__dfxtp_2 _5059_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[46][3] ),
    .D(_0054_));
 sky130_as_sc_hs__dfxtp_2 _5060_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[46][4] ),
    .D(_0055_));
 sky130_as_sc_hs__dfxtp_2 _5061_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[46][5] ),
    .D(_0056_));
 sky130_as_sc_hs__dfxtp_2 _5062_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[19][0] ),
    .D(_0057_));
 sky130_as_sc_hs__dfxtp_2 _5063_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[19][1] ),
    .D(_0058_));
 sky130_as_sc_hs__dfxtp_2 _5064_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[19][2] ),
    .D(_0059_));
 sky130_as_sc_hs__dfxtp_2 _5065_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[19][3] ),
    .D(_0060_));
 sky130_as_sc_hs__dfxtp_2 _5066_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[19][4] ),
    .D(_0061_));
 sky130_as_sc_hs__dfxtp_2 _5067_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[19][5] ),
    .D(_0062_));
 sky130_as_sc_hs__dfxtp_2 _5068_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[47][0] ),
    .D(_0063_));
 sky130_as_sc_hs__dfxtp_2 _5069_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[47][1] ),
    .D(_0064_));
 sky130_as_sc_hs__dfxtp_2 _5070_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[47][2] ),
    .D(_0065_));
 sky130_as_sc_hs__dfxtp_2 _5071_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[47][3] ),
    .D(_0066_));
 sky130_as_sc_hs__dfxtp_2 _5072_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[47][4] ),
    .D(_0067_));
 sky130_as_sc_hs__dfxtp_2 _5073_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_10_clk),
    .Q(\RAM[47][5] ),
    .D(_0068_));
 sky130_as_sc_hs__dfxtp_2 _5074_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[29][0] ),
    .D(_0069_));
 sky130_as_sc_hs__dfxtp_2 _5075_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[29][1] ),
    .D(_0070_));
 sky130_as_sc_hs__dfxtp_2 _5076_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[29][2] ),
    .D(_0071_));
 sky130_as_sc_hs__dfxtp_2 _5077_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[29][3] ),
    .D(_0072_));
 sky130_as_sc_hs__dfxtp_2 _5078_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[29][4] ),
    .D(_0073_));
 sky130_as_sc_hs__dfxtp_2 _5079_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[29][5] ),
    .D(_0074_));
 sky130_as_sc_hs__dfxtp_2 _5080_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[48][0] ),
    .D(_0075_));
 sky130_as_sc_hs__dfxtp_2 _5081_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[48][1] ),
    .D(_0076_));
 sky130_as_sc_hs__dfxtp_2 _5082_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[48][2] ),
    .D(_0077_));
 sky130_as_sc_hs__dfxtp_2 _5083_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[48][3] ),
    .D(_0078_));
 sky130_as_sc_hs__dfxtp_2 _5084_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[48][4] ),
    .D(_0079_));
 sky130_as_sc_hs__dfxtp_2 _5085_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[48][5] ),
    .D(_0080_));
 sky130_as_sc_hs__dfxtp_2 _5086_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[39][0] ),
    .D(_0081_));
 sky130_as_sc_hs__dfxtp_2 _5087_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[39][1] ),
    .D(_0082_));
 sky130_as_sc_hs__dfxtp_2 _5088_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[39][2] ),
    .D(_0083_));
 sky130_as_sc_hs__dfxtp_2 _5089_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[39][3] ),
    .D(_0084_));
 sky130_as_sc_hs__dfxtp_2 _5090_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[39][4] ),
    .D(_0085_));
 sky130_as_sc_hs__dfxtp_2 _5091_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[39][5] ),
    .D(_0086_));
 sky130_as_sc_hs__dfxtp_2 _5092_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_23_clk),
    .Q(\ROM_dest[0] ),
    .D(_0018_));
 sky130_as_sc_hs__dfxtp_2 _5093_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_23_clk),
    .Q(\ROM_dest[1] ),
    .D(_0019_));
 sky130_as_sc_hs__dfxtp_2 _5094_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_23_clk),
    .Q(\ROM_dest[2] ),
    .D(_0020_));
 sky130_as_sc_hs__dfxtp_2 _5095_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[57][0] ),
    .D(_0087_));
 sky130_as_sc_hs__dfxtp_2 _5096_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[57][1] ),
    .D(_0088_));
 sky130_as_sc_hs__dfxtp_2 _5097_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(\RAM[57][2] ),
    .D(_0089_));
 sky130_as_sc_hs__dfxtp_2 _5098_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[57][3] ),
    .D(_0090_));
 sky130_as_sc_hs__dfxtp_2 _5099_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[57][4] ),
    .D(_0091_));
 sky130_as_sc_hs__dfxtp_2 _5100_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[57][5] ),
    .D(_0092_));
 sky130_as_sc_hs__dfxtp_2 _5101_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[4][0] ),
    .D(_0093_));
 sky130_as_sc_hs__dfxtp_2 _5102_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[4][1] ),
    .D(_0094_));
 sky130_as_sc_hs__dfxtp_2 _5103_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[4][2] ),
    .D(_0095_));
 sky130_as_sc_hs__dfxtp_2 _5104_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[4][3] ),
    .D(_0096_));
 sky130_as_sc_hs__dfxtp_2 _5105_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[4][4] ),
    .D(_0097_));
 sky130_as_sc_hs__dfxtp_2 _5106_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[4][5] ),
    .D(_0098_));
 sky130_as_sc_hs__dfxtp_2 _5107_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[54][0] ),
    .D(_0099_));
 sky130_as_sc_hs__dfxtp_2 _5108_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[54][1] ),
    .D(_0100_));
 sky130_as_sc_hs__dfxtp_2 _5109_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[54][2] ),
    .D(_0101_));
 sky130_as_sc_hs__dfxtp_2 _5110_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[54][3] ),
    .D(_0102_));
 sky130_as_sc_hs__dfxtp_2 _5111_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[54][4] ),
    .D(_0103_));
 sky130_as_sc_hs__dfxtp_2 _5112_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[54][5] ),
    .D(_0104_));
 sky130_as_sc_hs__dfxtp_2 _5113_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[55][0] ),
    .D(_0105_));
 sky130_as_sc_hs__dfxtp_2 _5114_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[55][1] ),
    .D(_0106_));
 sky130_as_sc_hs__dfxtp_2 _5115_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[55][2] ),
    .D(_0107_));
 sky130_as_sc_hs__dfxtp_2 _5116_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[55][3] ),
    .D(_0108_));
 sky130_as_sc_hs__dfxtp_2 _5117_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[55][4] ),
    .D(_0109_));
 sky130_as_sc_hs__dfxtp_2 _5118_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[55][5] ),
    .D(_0110_));
 sky130_as_sc_hs__dfxtp_2 _5119_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[38][0] ),
    .D(_0111_));
 sky130_as_sc_hs__dfxtp_2 _5120_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[38][1] ),
    .D(_0112_));
 sky130_as_sc_hs__dfxtp_2 _5121_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[38][2] ),
    .D(_0113_));
 sky130_as_sc_hs__dfxtp_2 _5122_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[38][3] ),
    .D(_0114_));
 sky130_as_sc_hs__dfxtp_2 _5123_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[38][4] ),
    .D(_0115_));
 sky130_as_sc_hs__dfxtp_2 _5124_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[38][5] ),
    .D(_0116_));
 sky130_as_sc_hs__dfxtp_2 _5125_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[53][0] ),
    .D(_0117_));
 sky130_as_sc_hs__dfxtp_2 _5126_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[53][1] ),
    .D(_0118_));
 sky130_as_sc_hs__dfxtp_2 _5127_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[53][2] ),
    .D(_0119_));
 sky130_as_sc_hs__dfxtp_2 _5128_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[53][3] ),
    .D(_0120_));
 sky130_as_sc_hs__dfxtp_2 _5129_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[53][4] ),
    .D(_0121_));
 sky130_as_sc_hs__dfxtp_2 _5130_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[53][5] ),
    .D(_0122_));
 sky130_as_sc_hs__dfxtp_2 _5131_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\RAM[58][0] ),
    .D(_0123_));
 sky130_as_sc_hs__dfxtp_2 _5132_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[58][1] ),
    .D(_0124_));
 sky130_as_sc_hs__dfxtp_2 _5133_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[58][2] ),
    .D(_0125_));
 sky130_as_sc_hs__dfxtp_2 _5134_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\RAM[58][3] ),
    .D(_0126_));
 sky130_as_sc_hs__dfxtp_2 _5135_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\RAM[58][4] ),
    .D(_0127_));
 sky130_as_sc_hs__dfxtp_2 _5136_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\RAM[58][5] ),
    .D(_0128_));
 sky130_as_sc_hs__dfxtp_2 _5137_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[42][0] ),
    .D(_0129_));
 sky130_as_sc_hs__dfxtp_2 _5138_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[42][1] ),
    .D(_0130_));
 sky130_as_sc_hs__dfxtp_2 _5139_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[42][2] ),
    .D(_0131_));
 sky130_as_sc_hs__dfxtp_2 _5140_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[42][3] ),
    .D(_0132_));
 sky130_as_sc_hs__dfxtp_2 _5141_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[42][4] ),
    .D(_0133_));
 sky130_as_sc_hs__dfxtp_2 _5142_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[42][5] ),
    .D(_0134_));
 sky130_as_sc_hs__dfxtp_2 _5143_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[40][0] ),
    .D(_0135_));
 sky130_as_sc_hs__dfxtp_2 _5144_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[40][1] ),
    .D(_0136_));
 sky130_as_sc_hs__dfxtp_2 _5145_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[40][2] ),
    .D(_0137_));
 sky130_as_sc_hs__dfxtp_2 _5146_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[40][3] ),
    .D(_0138_));
 sky130_as_sc_hs__dfxtp_2 _5147_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[40][4] ),
    .D(_0139_));
 sky130_as_sc_hs__dfxtp_2 _5148_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[40][5] ),
    .D(_0140_));
 sky130_as_sc_hs__dfxtp_2 _5149_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\MAR[5] ),
    .D(_0005_));
 sky130_as_sc_hs__dfxtp_2 _5150_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[52][0] ),
    .D(_0141_));
 sky130_as_sc_hs__dfxtp_2 _5151_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[52][1] ),
    .D(_0142_));
 sky130_as_sc_hs__dfxtp_2 _5152_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[52][2] ),
    .D(_0143_));
 sky130_as_sc_hs__dfxtp_2 _5153_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[52][3] ),
    .D(_0144_));
 sky130_as_sc_hs__dfxtp_2 _5154_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[52][4] ),
    .D(_0145_));
 sky130_as_sc_hs__dfxtp_2 _5155_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[52][5] ),
    .D(_0146_));
 sky130_as_sc_hs__dfxtp_2 _5156_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[51][0] ),
    .D(_0147_));
 sky130_as_sc_hs__dfxtp_2 _5157_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[51][1] ),
    .D(_0148_));
 sky130_as_sc_hs__dfxtp_2 _5158_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[51][2] ),
    .D(_0149_));
 sky130_as_sc_hs__dfxtp_2 _5159_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[51][3] ),
    .D(_0150_));
 sky130_as_sc_hs__dfxtp_2 _5160_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_7_clk),
    .Q(\RAM[51][4] ),
    .D(_0151_));
 sky130_as_sc_hs__dfxtp_2 _5161_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[51][5] ),
    .D(_0152_));
 sky130_as_sc_hs__dfxtp_2 _5162_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_6_clk),
    .Q(\RAM[41][0] ),
    .D(_0153_));
 sky130_as_sc_hs__dfxtp_2 _5163_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[41][1] ),
    .D(_0154_));
 sky130_as_sc_hs__dfxtp_2 _5164_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[41][2] ),
    .D(_0155_));
 sky130_as_sc_hs__dfxtp_2 _5165_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[41][3] ),
    .D(_0156_));
 sky130_as_sc_hs__dfxtp_2 _5166_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[41][4] ),
    .D(_0157_));
 sky130_as_sc_hs__dfxtp_2 _5167_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[41][5] ),
    .D(_0158_));
 sky130_as_sc_hs__dfxtp_2 _5168_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[3][0] ),
    .D(_0159_));
 sky130_as_sc_hs__dfxtp_2 _5169_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[3][1] ),
    .D(_0160_));
 sky130_as_sc_hs__dfxtp_2 _5170_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[3][2] ),
    .D(_0161_));
 sky130_as_sc_hs__dfxtp_2 _5171_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[3][3] ),
    .D(_0162_));
 sky130_as_sc_hs__dfxtp_2 _5172_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[3][4] ),
    .D(_0163_));
 sky130_as_sc_hs__dfxtp_2 _5173_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[3][5] ),
    .D(_0164_));
 sky130_as_sc_hs__dfxtp_2 _5174_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\instr_cycle[0] ),
    .D(_0021_));
 sky130_as_sc_hs__dfxtp_4 _5175_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_23_clk),
    .Q(\instr_cycle[1] ),
    .D(_0022_));
 sky130_as_sc_hs__dfxtp_2 _5176_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\instr_cycle[2] ),
    .D(_0023_));
 sky130_as_sc_hs__dfxtp_2 _5177_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[21][0] ),
    .D(_0165_));
 sky130_as_sc_hs__dfxtp_2 _5178_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[21][1] ),
    .D(_0166_));
 sky130_as_sc_hs__dfxtp_2 _5179_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[21][2] ),
    .D(_0167_));
 sky130_as_sc_hs__dfxtp_2 _5180_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[21][3] ),
    .D(_0168_));
 sky130_as_sc_hs__dfxtp_2 _5181_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[21][4] ),
    .D(_0169_));
 sky130_as_sc_hs__dfxtp_2 _5182_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[21][5] ),
    .D(_0170_));
 sky130_as_sc_hs__dfxtp_2 _5183_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[50][0] ),
    .D(_0171_));
 sky130_as_sc_hs__dfxtp_2 _5184_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[50][1] ),
    .D(_0172_));
 sky130_as_sc_hs__dfxtp_2 _5185_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[50][2] ),
    .D(_0173_));
 sky130_as_sc_hs__dfxtp_2 _5186_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[50][3] ),
    .D(_0174_));
 sky130_as_sc_hs__dfxtp_2 _5187_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[50][4] ),
    .D(_0175_));
 sky130_as_sc_hs__dfxtp_2 _5188_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[50][5] ),
    .D(_0176_));
 sky130_as_sc_hs__dfxtp_2 _5189_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[14][0] ),
    .D(_0177_));
 sky130_as_sc_hs__dfxtp_2 _5190_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[14][1] ),
    .D(_0178_));
 sky130_as_sc_hs__dfxtp_2 _5191_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[14][2] ),
    .D(_0179_));
 sky130_as_sc_hs__dfxtp_2 _5192_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[14][3] ),
    .D(_0180_));
 sky130_as_sc_hs__dfxtp_2 _5193_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[14][4] ),
    .D(_0181_));
 sky130_as_sc_hs__dfxtp_2 _5194_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[14][5] ),
    .D(_0182_));
 sky130_as_sc_hs__dfxtp_2 _5195_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[37][0] ),
    .D(_0183_));
 sky130_as_sc_hs__dfxtp_2 _5196_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[37][1] ),
    .D(_0184_));
 sky130_as_sc_hs__dfxtp_2 _5197_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[37][2] ),
    .D(_0185_));
 sky130_as_sc_hs__dfxtp_2 _5198_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[37][3] ),
    .D(_0186_));
 sky130_as_sc_hs__dfxtp_2 _5199_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[37][4] ),
    .D(_0187_));
 sky130_as_sc_hs__dfxtp_2 _5200_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[37][5] ),
    .D(_0188_));
 sky130_as_sc_hs__dfxtp_2 _5201_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[15][0] ),
    .D(_0189_));
 sky130_as_sc_hs__dfxtp_2 _5202_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\RAM[15][1] ),
    .D(_0190_));
 sky130_as_sc_hs__dfxtp_2 _5203_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[15][2] ),
    .D(_0191_));
 sky130_as_sc_hs__dfxtp_2 _5204_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[15][3] ),
    .D(_0192_));
 sky130_as_sc_hs__dfxtp_2 _5205_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\RAM[15][4] ),
    .D(_0193_));
 sky130_as_sc_hs__dfxtp_2 _5206_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[15][5] ),
    .D(_0194_));
 sky130_as_sc_hs__dfxtp_2 _5207_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[36][0] ),
    .D(_0195_));
 sky130_as_sc_hs__dfxtp_2 _5208_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[36][1] ),
    .D(_0196_));
 sky130_as_sc_hs__dfxtp_2 _5209_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[36][2] ),
    .D(_0197_));
 sky130_as_sc_hs__dfxtp_2 _5210_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_3_clk),
    .Q(\RAM[36][3] ),
    .D(_0198_));
 sky130_as_sc_hs__dfxtp_2 _5211_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[36][4] ),
    .D(_0199_));
 sky130_as_sc_hs__dfxtp_2 _5212_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[36][5] ),
    .D(_0200_));
 sky130_as_sc_hs__dfxtp_2 _5213_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[16][0] ),
    .D(_0201_));
 sky130_as_sc_hs__dfxtp_2 _5214_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[16][1] ),
    .D(_0202_));
 sky130_as_sc_hs__dfxtp_2 _5215_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[16][2] ),
    .D(_0203_));
 sky130_as_sc_hs__dfxtp_2 _5216_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[16][3] ),
    .D(_0204_));
 sky130_as_sc_hs__dfxtp_2 _5217_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[16][4] ),
    .D(_0205_));
 sky130_as_sc_hs__dfxtp_2 _5218_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[16][5] ),
    .D(_0206_));
 sky130_as_sc_hs__dfxtp_2 _5219_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[35][0] ),
    .D(_0207_));
 sky130_as_sc_hs__dfxtp_2 _5220_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[35][1] ),
    .D(_0208_));
 sky130_as_sc_hs__dfxtp_2 _5221_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[35][2] ),
    .D(_0209_));
 sky130_as_sc_hs__dfxtp_2 _5222_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[35][3] ),
    .D(_0210_));
 sky130_as_sc_hs__dfxtp_2 _5223_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[35][4] ),
    .D(_0211_));
 sky130_as_sc_hs__dfxtp_2 _5224_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[35][5] ),
    .D(_0212_));
 sky130_as_sc_hs__dfxtp_2 _5225_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_2_clk),
    .Q(\RAM[17][0] ),
    .D(_0213_));
 sky130_as_sc_hs__dfxtp_2 _5226_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[17][1] ),
    .D(_0214_));
 sky130_as_sc_hs__dfxtp_2 _5227_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[17][2] ),
    .D(_0215_));
 sky130_as_sc_hs__dfxtp_2 _5228_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[17][3] ),
    .D(_0216_));
 sky130_as_sc_hs__dfxtp_2 _5229_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[17][4] ),
    .D(_0217_));
 sky130_as_sc_hs__dfxtp_2 _5230_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[17][5] ),
    .D(_0218_));
 sky130_as_sc_hs__dfxtp_2 _5231_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[34][0] ),
    .D(_0219_));
 sky130_as_sc_hs__dfxtp_2 _5232_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[34][1] ),
    .D(_0220_));
 sky130_as_sc_hs__dfxtp_2 _5233_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[34][2] ),
    .D(_0221_));
 sky130_as_sc_hs__dfxtp_2 _5234_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[34][3] ),
    .D(_0222_));
 sky130_as_sc_hs__dfxtp_2 _5235_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[34][4] ),
    .D(_0223_));
 sky130_as_sc_hs__dfxtp_2 _5236_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[34][5] ),
    .D(_0224_));
 sky130_as_sc_hs__dfxtp_2 _5237_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[18][0] ),
    .D(_0225_));
 sky130_as_sc_hs__dfxtp_2 _5238_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[18][1] ),
    .D(_0226_));
 sky130_as_sc_hs__dfxtp_2 _5239_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[18][2] ),
    .D(_0227_));
 sky130_as_sc_hs__dfxtp_2 _5240_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_1_clk),
    .Q(\RAM[18][3] ),
    .D(_0228_));
 sky130_as_sc_hs__dfxtp_2 _5241_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[18][4] ),
    .D(_0229_));
 sky130_as_sc_hs__dfxtp_2 _5242_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[18][5] ),
    .D(_0230_));
 sky130_as_sc_hs__dfxtp_2 _5243_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[33][0] ),
    .D(_0231_));
 sky130_as_sc_hs__dfxtp_2 _5244_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[33][1] ),
    .D(_0232_));
 sky130_as_sc_hs__dfxtp_2 _5245_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[33][2] ),
    .D(_0233_));
 sky130_as_sc_hs__dfxtp_2 _5246_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[33][3] ),
    .D(_0234_));
 sky130_as_sc_hs__dfxtp_2 _5247_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[33][4] ),
    .D(_0235_));
 sky130_as_sc_hs__dfxtp_2 _5248_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[33][5] ),
    .D(_0236_));
 sky130_as_sc_hs__dfxtp_2 _5249_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[1][0] ),
    .D(_0237_));
 sky130_as_sc_hs__dfxtp_2 _5250_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[1][1] ),
    .D(_0238_));
 sky130_as_sc_hs__dfxtp_2 _5251_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[1][2] ),
    .D(_0239_));
 sky130_as_sc_hs__dfxtp_2 _5252_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[1][3] ),
    .D(_0240_));
 sky130_as_sc_hs__dfxtp_2 _5253_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[1][4] ),
    .D(_0241_));
 sky130_as_sc_hs__dfxtp_2 _5254_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[1][5] ),
    .D(_0242_));
 sky130_as_sc_hs__dfxtp_2 _5255_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[32][0] ),
    .D(_0243_));
 sky130_as_sc_hs__dfxtp_2 _5256_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[32][1] ),
    .D(_0244_));
 sky130_as_sc_hs__dfxtp_2 _5257_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[32][2] ),
    .D(_0245_));
 sky130_as_sc_hs__dfxtp_2 _5258_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[32][3] ),
    .D(_0246_));
 sky130_as_sc_hs__dfxtp_2 _5259_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[32][4] ),
    .D(_0247_));
 sky130_as_sc_hs__dfxtp_2 _5260_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_36_clk),
    .Q(\RAM[32][5] ),
    .D(_0248_));
 sky130_as_sc_hs__dfxtp_2 _5261_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[20][0] ),
    .D(_0249_));
 sky130_as_sc_hs__dfxtp_2 _5262_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[20][1] ),
    .D(_0250_));
 sky130_as_sc_hs__dfxtp_2 _5263_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[20][2] ),
    .D(_0251_));
 sky130_as_sc_hs__dfxtp_2 _5264_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[20][3] ),
    .D(_0252_));
 sky130_as_sc_hs__dfxtp_2 _5265_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[20][4] ),
    .D(_0253_));
 sky130_as_sc_hs__dfxtp_2 _5266_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[20][5] ),
    .D(_0254_));
 sky130_as_sc_hs__dfxtp_2 _5267_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[31][0] ),
    .D(_0255_));
 sky130_as_sc_hs__dfxtp_2 _5268_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[31][1] ),
    .D(_0256_));
 sky130_as_sc_hs__dfxtp_2 _5269_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[31][2] ),
    .D(_0257_));
 sky130_as_sc_hs__dfxtp_2 _5270_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[31][3] ),
    .D(_0258_));
 sky130_as_sc_hs__dfxtp_2 _5271_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[31][4] ),
    .D(_0259_));
 sky130_as_sc_hs__dfxtp_2 _5272_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[31][5] ),
    .D(_0260_));
 sky130_as_sc_hs__dfxtp_2 _5273_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[30][0] ),
    .D(_0261_));
 sky130_as_sc_hs__dfxtp_2 _5274_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[30][1] ),
    .D(_0262_));
 sky130_as_sc_hs__dfxtp_2 _5275_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[30][2] ),
    .D(_0263_));
 sky130_as_sc_hs__dfxtp_2 _5276_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[30][3] ),
    .D(_0264_));
 sky130_as_sc_hs__dfxtp_2 _5277_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[30][4] ),
    .D(_0265_));
 sky130_as_sc_hs__dfxtp_2 _5278_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[30][5] ),
    .D(_0266_));
 sky130_as_sc_hs__dfxtp_4 _5279_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(uio_out[0]),
    .D(_0267_));
 sky130_as_sc_hs__dfxtp_4 _5280_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uio_out[1]),
    .D(_0268_));
 sky130_as_sc_hs__dfxtp_4 _5281_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uio_out[2]),
    .D(_0269_));
 sky130_as_sc_hs__dfxtp_4 _5282_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uio_out[3]),
    .D(_0270_));
 sky130_as_sc_hs__dfxtp_4 _5283_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uio_out[4]),
    .D(_0271_));
 sky130_as_sc_hs__dfxtp_4 _5284_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uio_out[5]),
    .D(_0272_));
 sky130_as_sc_hs__dfxtp_2 _5285_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[2][0] ),
    .D(_0273_));
 sky130_as_sc_hs__dfxtp_2 _5286_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[2][1] ),
    .D(_0274_));
 sky130_as_sc_hs__dfxtp_2 _5287_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[2][2] ),
    .D(_0275_));
 sky130_as_sc_hs__dfxtp_2 _5288_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[2][3] ),
    .D(_0276_));
 sky130_as_sc_hs__dfxtp_2 _5289_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[2][4] ),
    .D(_0277_));
 sky130_as_sc_hs__dfxtp_2 _5290_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[2][5] ),
    .D(_0278_));
 sky130_as_sc_hs__dfxtp_2 _5291_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[6][0] ),
    .D(_0279_));
 sky130_as_sc_hs__dfxtp_2 _5292_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[6][1] ),
    .D(_0280_));
 sky130_as_sc_hs__dfxtp_2 _5293_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[6][2] ),
    .D(_0281_));
 sky130_as_sc_hs__dfxtp_2 _5294_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[6][3] ),
    .D(_0282_));
 sky130_as_sc_hs__dfxtp_2 _5295_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[6][4] ),
    .D(_0283_));
 sky130_as_sc_hs__dfxtp_2 _5296_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[6][5] ),
    .D(_0284_));
 sky130_as_sc_hs__dfxtp_2 _5297_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[28][0] ),
    .D(_0285_));
 sky130_as_sc_hs__dfxtp_2 _5298_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[28][1] ),
    .D(_0286_));
 sky130_as_sc_hs__dfxtp_2 _5299_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[28][2] ),
    .D(_0287_));
 sky130_as_sc_hs__dfxtp_2 _5300_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[28][3] ),
    .D(_0288_));
 sky130_as_sc_hs__dfxtp_2 _5301_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[28][4] ),
    .D(_0289_));
 sky130_as_sc_hs__dfxtp_2 _5302_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[28][5] ),
    .D(_0290_));
 sky130_as_sc_hs__dfxtp_2 _5303_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[7][0] ),
    .D(_0291_));
 sky130_as_sc_hs__dfxtp_2 _5304_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[7][1] ),
    .D(_0292_));
 sky130_as_sc_hs__dfxtp_2 _5305_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[7][2] ),
    .D(_0293_));
 sky130_as_sc_hs__dfxtp_2 _5306_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[7][3] ),
    .D(_0294_));
 sky130_as_sc_hs__dfxtp_2 _5307_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_33_clk),
    .Q(\RAM[7][4] ),
    .D(_0295_));
 sky130_as_sc_hs__dfxtp_2 _5308_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[7][5] ),
    .D(_0296_));
 sky130_as_sc_hs__dfxtp_2 _5309_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[27][0] ),
    .D(_0297_));
 sky130_as_sc_hs__dfxtp_2 _5310_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[27][1] ),
    .D(_0298_));
 sky130_as_sc_hs__dfxtp_2 _5311_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[27][2] ),
    .D(_0299_));
 sky130_as_sc_hs__dfxtp_2 _5312_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[27][3] ),
    .D(_0300_));
 sky130_as_sc_hs__dfxtp_2 _5313_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[27][4] ),
    .D(_0301_));
 sky130_as_sc_hs__dfxtp_2 _5314_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[27][5] ),
    .D(_0302_));
 sky130_as_sc_hs__dfxtp_2 _5315_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[8][0] ),
    .D(_0303_));
 sky130_as_sc_hs__dfxtp_2 _5316_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[8][1] ),
    .D(_0304_));
 sky130_as_sc_hs__dfxtp_2 _5317_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[8][2] ),
    .D(_0305_));
 sky130_as_sc_hs__dfxtp_2 _5318_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[8][3] ),
    .D(_0306_));
 sky130_as_sc_hs__dfxtp_2 _5319_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[8][4] ),
    .D(_0307_));
 sky130_as_sc_hs__dfxtp_2 _5320_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[8][5] ),
    .D(_0308_));
 sky130_as_sc_hs__dfxtp_2 _5321_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[26][0] ),
    .D(_0309_));
 sky130_as_sc_hs__dfxtp_2 _5322_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[26][1] ),
    .D(_0310_));
 sky130_as_sc_hs__dfxtp_2 _5323_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[26][2] ),
    .D(_0311_));
 sky130_as_sc_hs__dfxtp_2 _5324_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[26][3] ),
    .D(_0312_));
 sky130_as_sc_hs__dfxtp_2 _5325_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[26][4] ),
    .D(_0313_));
 sky130_as_sc_hs__dfxtp_2 _5326_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[26][5] ),
    .D(_0314_));
 sky130_as_sc_hs__dfxtp_4 _5327_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(uio_oe[0]),
    .D(_0315_));
 sky130_as_sc_hs__dfxtp_4 _5328_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(uio_oe[1]),
    .D(_0316_));
 sky130_as_sc_hs__dfxtp_4 _5329_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uio_oe[2]),
    .D(_0317_));
 sky130_as_sc_hs__dfxtp_4 _5330_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(uio_oe[3]),
    .D(_0318_));
 sky130_as_sc_hs__dfxtp_4 _5331_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uio_oe[4]),
    .D(_0319_));
 sky130_as_sc_hs__dfxtp_4 _5332_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(uio_oe[5]),
    .D(_0320_));
 sky130_as_sc_hs__dfxtp_2 _5333_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[0][0] ),
    .D(_0321_));
 sky130_as_sc_hs__dfxtp_2 _5334_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[0][1] ),
    .D(_0322_));
 sky130_as_sc_hs__dfxtp_2 _5335_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_0_clk),
    .Q(\RAM[0][2] ),
    .D(_0323_));
 sky130_as_sc_hs__dfxtp_2 _5336_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[0][3] ),
    .D(_0324_));
 sky130_as_sc_hs__dfxtp_2 _5337_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_35_clk),
    .Q(\RAM[0][4] ),
    .D(_0325_));
 sky130_as_sc_hs__dfxtp_2 _5338_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_34_clk),
    .Q(\RAM[0][5] ),
    .D(_0326_));
 sky130_as_sc_hs__dfxtp_2 _5339_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[25][0] ),
    .D(_0327_));
 sky130_as_sc_hs__dfxtp_2 _5340_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[25][1] ),
    .D(_0328_));
 sky130_as_sc_hs__dfxtp_2 _5341_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[25][2] ),
    .D(_0329_));
 sky130_as_sc_hs__dfxtp_2 _5342_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[25][3] ),
    .D(_0330_));
 sky130_as_sc_hs__dfxtp_2 _5343_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[25][4] ),
    .D(_0331_));
 sky130_as_sc_hs__dfxtp_2 _5344_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[25][5] ),
    .D(_0332_));
 sky130_as_sc_hs__dfxtp_4 _5345_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(uo_out[0]),
    .D(_0333_));
 sky130_as_sc_hs__dfxtp_4 _5346_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(uo_out[1]),
    .D(_0334_));
 sky130_as_sc_hs__dfxtp_4 _5347_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uo_out[2]),
    .D(_0335_));
 sky130_as_sc_hs__dfxtp_4 _5348_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uo_out[3]),
    .D(_0336_));
 sky130_as_sc_hs__dfxtp_4 _5349_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uo_out[4]),
    .D(_0337_));
 sky130_as_sc_hs__dfxtp_4 _5350_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(uo_out[5]),
    .D(_0338_));
 sky130_as_sc_hs__dfxtp_2 _5351_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[10][0] ),
    .D(_0339_));
 sky130_as_sc_hs__dfxtp_2 _5352_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[10][1] ),
    .D(_0340_));
 sky130_as_sc_hs__dfxtp_2 _5353_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[10][2] ),
    .D(_0341_));
 sky130_as_sc_hs__dfxtp_2 _5354_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[10][3] ),
    .D(_0342_));
 sky130_as_sc_hs__dfxtp_2 _5355_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[10][4] ),
    .D(_0343_));
 sky130_as_sc_hs__dfxtp_2 _5356_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[10][5] ),
    .D(_0344_));
 sky130_as_sc_hs__dfxtp_2 _5357_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_15_clk),
    .Q(\RAM[56][0] ),
    .D(_0345_));
 sky130_as_sc_hs__dfxtp_2 _5358_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_15_clk),
    .Q(\RAM[56][1] ),
    .D(_0346_));
 sky130_as_sc_hs__dfxtp_2 _5359_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\RAM[56][2] ),
    .D(_0347_));
 sky130_as_sc_hs__dfxtp_2 _5360_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_15_clk),
    .Q(\RAM[56][3] ),
    .D(_0348_));
 sky130_as_sc_hs__dfxtp_2 _5361_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\RAM[56][4] ),
    .D(_0349_));
 sky130_as_sc_hs__dfxtp_2 _5362_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\RAM[56][5] ),
    .D(_0350_));
 sky130_as_sc_hs__dfxtp_2 _5363_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[5][0] ),
    .D(_0351_));
 sky130_as_sc_hs__dfxtp_2 _5364_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[5][1] ),
    .D(_0352_));
 sky130_as_sc_hs__dfxtp_2 _5365_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[5][2] ),
    .D(_0353_));
 sky130_as_sc_hs__dfxtp_2 _5366_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[5][3] ),
    .D(_0354_));
 sky130_as_sc_hs__dfxtp_2 _5367_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[5][4] ),
    .D(_0355_));
 sky130_as_sc_hs__dfxtp_2 _5368_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[5][5] ),
    .D(_0356_));
 sky130_as_sc_hs__dfxtp_2 _5369_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[24][0] ),
    .D(_0357_));
 sky130_as_sc_hs__dfxtp_2 _5370_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[24][1] ),
    .D(_0358_));
 sky130_as_sc_hs__dfxtp_2 _5371_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[24][2] ),
    .D(_0359_));
 sky130_as_sc_hs__dfxtp_2 _5372_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_29_clk),
    .Q(\RAM[24][3] ),
    .D(_0360_));
 sky130_as_sc_hs__dfxtp_2 _5373_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[24][4] ),
    .D(_0361_));
 sky130_as_sc_hs__dfxtp_2 _5374_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_28_clk),
    .Q(\RAM[24][5] ),
    .D(_0362_));
 sky130_as_sc_hs__dfxtp_2 _5375_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[11][0] ),
    .D(_0363_));
 sky130_as_sc_hs__dfxtp_2 _5376_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\RAM[11][1] ),
    .D(_0364_));
 sky130_as_sc_hs__dfxtp_2 _5377_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[11][2] ),
    .D(_0365_));
 sky130_as_sc_hs__dfxtp_2 _5378_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[11][3] ),
    .D(_0366_));
 sky130_as_sc_hs__dfxtp_2 _5379_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[11][4] ),
    .D(_0367_));
 sky130_as_sc_hs__dfxtp_2 _5380_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[11][5] ),
    .D(_0368_));
 sky130_as_sc_hs__dfxtp_2 _5381_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[23][0] ),
    .D(_0369_));
 sky130_as_sc_hs__dfxtp_2 _5382_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[23][1] ),
    .D(_0370_));
 sky130_as_sc_hs__dfxtp_2 _5383_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[23][2] ),
    .D(_0371_));
 sky130_as_sc_hs__dfxtp_2 _5384_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[23][3] ),
    .D(_0372_));
 sky130_as_sc_hs__dfxtp_2 _5385_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[23][4] ),
    .D(_0373_));
 sky130_as_sc_hs__dfxtp_2 _5386_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_32_clk),
    .Q(\RAM[23][5] ),
    .D(_0374_));
 sky130_as_sc_hs__dfxtp_2 _5387_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[12][0] ),
    .D(_0375_));
 sky130_as_sc_hs__dfxtp_2 _5388_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[12][1] ),
    .D(_0376_));
 sky130_as_sc_hs__dfxtp_2 _5389_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[12][2] ),
    .D(_0377_));
 sky130_as_sc_hs__dfxtp_2 _5390_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[12][3] ),
    .D(_0378_));
 sky130_as_sc_hs__dfxtp_2 _5391_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[12][4] ),
    .D(_0379_));
 sky130_as_sc_hs__dfxtp_2 _5392_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[12][5] ),
    .D(_0380_));
 sky130_as_sc_hs__dfxtp_2 _5393_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[22][0] ),
    .D(_0381_));
 sky130_as_sc_hs__dfxtp_2 _5394_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[22][1] ),
    .D(_0382_));
 sky130_as_sc_hs__dfxtp_2 _5395_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[22][2] ),
    .D(_0383_));
 sky130_as_sc_hs__dfxtp_2 _5396_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_5_clk),
    .Q(\RAM[22][3] ),
    .D(_0384_));
 sky130_as_sc_hs__dfxtp_2 _5397_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[22][4] ),
    .D(_0385_));
 sky130_as_sc_hs__dfxtp_2 _5398_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_4_clk),
    .Q(\RAM[22][5] ),
    .D(_0386_));
 sky130_as_sc_hs__dfxtp_2 _5399_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[13][0] ),
    .D(_0387_));
 sky130_as_sc_hs__dfxtp_2 _5400_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\RAM[13][1] ),
    .D(_0388_));
 sky130_as_sc_hs__dfxtp_2 _5401_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[13][2] ),
    .D(_0389_));
 sky130_as_sc_hs__dfxtp_2 _5402_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[13][3] ),
    .D(_0390_));
 sky130_as_sc_hs__dfxtp_2 _5403_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\RAM[13][4] ),
    .D(_0391_));
 sky130_as_sc_hs__dfxtp_2 _5404_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_30_clk),
    .Q(\RAM[13][5] ),
    .D(_0392_));
 sky130_as_sc_hs__dfxtp_2 _5405_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(\RAM[61][0] ),
    .D(_0393_));
 sky130_as_sc_hs__dfxtp_2 _5406_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[61][1] ),
    .D(_0394_));
 sky130_as_sc_hs__dfxtp_2 _5407_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(\RAM[61][2] ),
    .D(_0395_));
 sky130_as_sc_hs__dfxtp_2 _5408_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(\RAM[61][3] ),
    .D(_0396_));
 sky130_as_sc_hs__dfxtp_2 _5409_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(\RAM[61][4] ),
    .D(_0397_));
 sky130_as_sc_hs__dfxtp_2 _5410_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_11_clk),
    .Q(\RAM[61][5] ),
    .D(_0398_));
 sky130_as_sc_hs__dfxtp_2 _5411_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\A[0] ),
    .D(_0399_));
 sky130_as_sc_hs__dfxtp_2 _5412_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\A[1] ),
    .D(_0400_));
 sky130_as_sc_hs__dfxtp_2 _5413_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\A[2] ),
    .D(_0401_));
 sky130_as_sc_hs__dfxtp_4 _5414_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\A[3] ),
    .D(_0402_));
 sky130_as_sc_hs__dfxtp_2 _5415_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\A[4] ),
    .D(_0403_));
 sky130_as_sc_hs__dfxtp_2 _5416_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\A[5] ),
    .D(_0404_));
 sky130_as_sc_hs__dfxtp_2 _5417_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\B[0] ),
    .D(_0405_));
 sky130_as_sc_hs__dfxtp_2 _5418_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\B[1] ),
    .D(_0406_));
 sky130_as_sc_hs__dfxtp_2 _5419_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\B[2] ),
    .D(_0407_));
 sky130_as_sc_hs__dfxtp_2 _5420_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\B[3] ),
    .D(_0408_));
 sky130_as_sc_hs__dfxtp_2 _5421_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\B[4] ),
    .D(_0409_));
 sky130_as_sc_hs__dfxtp_2 _5422_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\B[5] ),
    .D(_0410_));
 sky130_as_sc_hs__dfxtp_2 _5423_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\P[0] ),
    .D(_0006_));
 sky130_as_sc_hs__dfxtp_2 _5424_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\P[1] ),
    .D(_0007_));
 sky130_as_sc_hs__dfxtp_2 _5425_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\P[2] ),
    .D(_0008_));
 sky130_as_sc_hs__dfxtp_2 _5426_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\P[3] ),
    .D(_0009_));
 sky130_as_sc_hs__dfxtp_2 _5427_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\P[4] ),
    .D(_0010_));
 sky130_as_sc_hs__dfxtp_2 _5428_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\P[5] ),
    .D(_0011_));
 sky130_as_sc_hs__dfxtp_4 _5429_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_24_clk),
    .Q(carry),
    .D(_0411_));
 sky130_as_sc_hs__dfxtp_4 _5430_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_24_clk),
    .Q(zero),
    .D(_0412_));
 sky130_as_sc_hs__dfxtp_2 _5431_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\MAR[0] ),
    .D(_0000_));
 sky130_as_sc_hs__dfxtp_2 _5432_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\MAR[1] ),
    .D(_0001_));
 sky130_as_sc_hs__dfxtp_2 _5433_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\MAR[2] ),
    .D(_0002_));
 sky130_as_sc_hs__dfxtp_2 _5434_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\MAR[3] ),
    .D(_0003_));
 sky130_as_sc_hs__dfxtp_2 _5435_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\MAR[4] ),
    .D(_0004_));
 sky130_as_sc_hs__dfxtp_2 _5436_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\PC[0] ),
    .D(_0413_));
 sky130_as_sc_hs__dfxtp_2 _5437_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\PC[1] ),
    .D(_0414_));
 sky130_as_sc_hs__dfxtp_4 _5438_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_23_clk),
    .Q(\PC[2] ),
    .D(_0415_));
 sky130_as_sc_hs__dfxtp_2 _5439_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\PC[3] ),
    .D(_0416_));
 sky130_as_sc_hs__dfxtp_4 _5440_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\PC[4] ),
    .D(_0417_));
 sky130_as_sc_hs__dfxtp_4 _5441_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\PC[5] ),
    .D(_0418_));
 sky130_as_sc_hs__dfxtp_2 _5442_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\PC[6] ),
    .D(_0419_));
 sky130_as_sc_hs__dfxtp_2 _5443_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\PC[7] ),
    .D(_0420_));
 sky130_as_sc_hs__dfxtp_2 _5444_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\PC[8] ),
    .D(_0421_));
 sky130_as_sc_hs__dfxtp_2 _5445_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\PC[9] ),
    .D(_0422_));
 sky130_as_sc_hs__dfxtp_2 _5446_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\PC[10] ),
    .D(_0423_));
 sky130_as_sc_hs__dfxtp_2 _5447_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\PC[11] ),
    .D(_0424_));
 sky130_as_sc_hs__dfxtp_2 _5448_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\insin[0] ),
    .D(_0012_));
 sky130_as_sc_hs__dfxtp_2 _5449_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\insin[1] ),
    .D(_0013_));
 sky130_as_sc_hs__dfxtp_2 _5450_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\insin[2] ),
    .D(_0014_));
 sky130_as_sc_hs__dfxtp_2 _5451_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\insin[3] ),
    .D(_0015_));
 sky130_as_sc_hs__dfxtp_2 _5452_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\insin[4] ),
    .D(_0016_));
 sky130_as_sc_hs__dfxtp_2 _5453_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_17_clk),
    .Q(\insin[5] ),
    .D(_0017_));
 sky130_as_sc_hs__dfxtp_2 _5454_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_24_clk),
    .Q(compat),
    .D(_0425_));
 sky130_as_sc_hs__dfxtp_2 _5455_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\imm_buff[0] ),
    .D(_0426_));
 sky130_as_sc_hs__dfxtp_2 _5456_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\imm_buff[1] ),
    .D(_0427_));
 sky130_as_sc_hs__dfxtp_2 _5457_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_15_clk),
    .Q(\imm_buff[2] ),
    .D(_0428_));
 sky130_as_sc_hs__dfxtp_2 _5458_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\imm_buff[3] ),
    .D(_0429_));
 sky130_as_sc_hs__dfxtp_2 _5459_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_15_clk),
    .Q(\imm_buff[4] ),
    .D(_0430_));
 sky130_as_sc_hs__dfxtp_2 _5460_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\imm_buff[5] ),
    .D(_0431_));
 sky130_as_sc_hs__dfxtp_2 _5461_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\last_PC[0] ),
    .D(_0432_));
 sky130_as_sc_hs__dfxtp_2 _5462_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\last_PC[1] ),
    .D(_0433_));
 sky130_as_sc_hs__dfxtp_2 _5463_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_24_clk),
    .Q(\last_PC[2] ),
    .D(_0434_));
 sky130_as_sc_hs__dfxtp_2 _5464_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\last_PC[3] ),
    .D(_0435_));
 sky130_as_sc_hs__dfxtp_2 _5465_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\last_PC[4] ),
    .D(_0436_));
 sky130_as_sc_hs__dfxtp_2 _5466_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\last_PC[5] ),
    .D(_0437_));
 sky130_as_sc_hs__dfxtp_2 _5467_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\last_PC[6] ),
    .D(_0438_));
 sky130_as_sc_hs__dfxtp_2 _5468_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_22_clk),
    .Q(\last_PC[7] ),
    .D(_0439_));
 sky130_as_sc_hs__dfxtp_2 _5469_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\last_PC[8] ),
    .D(_0440_));
 sky130_as_sc_hs__dfxtp_2 _5470_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\last_PC[9] ),
    .D(_0441_));
 sky130_as_sc_hs__dfxtp_2 _5471_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\last_PC[10] ),
    .D(_0442_));
 sky130_as_sc_hs__dfxtp_2 _5472_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_23_clk),
    .Q(\last_PC[11] ),
    .D(_0443_));
 sky130_as_sc_hs__dfxtp_2 _5473_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_24_clk),
    .Q(\last_flags[0] ),
    .D(_0444_));
 sky130_as_sc_hs__dfxtp_2 _5474_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_24_clk),
    .Q(\last_flags[1] ),
    .D(_0445_));
 sky130_as_sc_hs__dfxtp_2 _5475_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\last_A[0] ),
    .D(_0446_));
 sky130_as_sc_hs__dfxtp_2 _5476_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_25_clk),
    .Q(\last_A[1] ),
    .D(_0447_));
 sky130_as_sc_hs__dfxtp_2 _5477_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\last_A[2] ),
    .D(_0448_));
 sky130_as_sc_hs__dfxtp_2 _5478_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\last_A[3] ),
    .D(_0449_));
 sky130_as_sc_hs__dfxtp_2 _5479_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\last_A[4] ),
    .D(_0450_));
 sky130_as_sc_hs__dfxtp_2 _5480_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\last_A[5] ),
    .D(_0451_));
 sky130_as_sc_hs__dfxtp_2 _5481_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\last_B[0] ),
    .D(_0452_));
 sky130_as_sc_hs__dfxtp_2 _5482_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\last_B[1] ),
    .D(_0453_));
 sky130_as_sc_hs__dfxtp_2 _5483_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\last_B[2] ),
    .D(_0454_));
 sky130_as_sc_hs__dfxtp_2 _5484_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\last_B[3] ),
    .D(_0455_));
 sky130_as_sc_hs__dfxtp_2 _5485_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\last_B[4] ),
    .D(_0456_));
 sky130_as_sc_hs__dfxtp_2 _5486_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\last_B[5] ),
    .D(_0457_));
 sky130_as_sc_hs__dfxtp_2 _5487_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\last_MAR[0] ),
    .D(_0458_));
 sky130_as_sc_hs__dfxtp_2 _5488_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_16_clk),
    .Q(\last_MAR[1] ),
    .D(_0459_));
 sky130_as_sc_hs__dfxtp_2 _5489_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_17_clk),
    .Q(\last_MAR[2] ),
    .D(_0460_));
 sky130_as_sc_hs__dfxtp_2 _5490_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_15_clk),
    .Q(\last_MAR[3] ),
    .D(_0461_));
 sky130_as_sc_hs__dfxtp_2 _5491_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_15_clk),
    .Q(\last_MAR[4] ),
    .D(_0462_));
 sky130_as_sc_hs__dfxtp_2 _5492_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_17_clk),
    .Q(\last_MAR[5] ),
    .D(_0463_));
 sky130_as_sc_hs__dfxtp_2 _5493_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\last_P[0] ),
    .D(_0464_));
 sky130_as_sc_hs__dfxtp_2 _5494_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\last_P[1] ),
    .D(_0465_));
 sky130_as_sc_hs__dfxtp_2 _5495_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_17_clk),
    .Q(\last_P[2] ),
    .D(_0466_));
 sky130_as_sc_hs__dfxtp_2 _5496_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\last_P[3] ),
    .D(_0467_));
 sky130_as_sc_hs__dfxtp_2 _5497_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_17_clk),
    .Q(\last_P[4] ),
    .D(_0468_));
 sky130_as_sc_hs__dfxtp_2 _5498_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_17_clk),
    .Q(\last_P[5] ),
    .D(_0469_));
 sky130_as_sc_hs__dfxtp_2 _5499_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_17_clk),
    .Q(needs_irupt),
    .D(_0470_));
 sky130_as_sc_hs__dfxtp_2 _5500_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_23_clk),
    .Q(in_irupt),
    .D(_0471_));
 sky130_as_sc_hs__dfxtp_4 _5501_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(\ROM_spi_cycle[0] ),
    .D(_0472_));
 sky130_as_sc_hs__dfxtp_2 _5502_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(\ROM_spi_cycle[1] ),
    .D(_0473_));
 sky130_as_sc_hs__dfxtp_2 _5503_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(\ROM_spi_cycle[2] ),
    .D(_0474_));
 sky130_as_sc_hs__dfxtp_2 _5504_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(\ROM_spi_cycle[3] ),
    .D(_0475_));
 sky130_as_sc_hs__dfxtp_2 _5505_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(\ROM_spi_cycle[4] ),
    .D(_0476_));
 sky130_as_sc_hs__dfxtp_2 _5506_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(last_inter),
    .D(_0477_));
 sky130_as_sc_hs__dfxtp_2 _5507_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(CS_ROM),
    .D(_0478_));
 sky130_as_sc_hs__dfxtp_2 _5508_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(SCLK_ROM),
    .D(_0479_));
 sky130_as_sc_hs__dfxtp_2 _5509_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(ROM_DO),
    .D(_0480_));
 sky130_as_sc_hs__dfxtp_2 _5510_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\ROM_spi_dat_out[0] ),
    .D(_0481_));
 sky130_as_sc_hs__dfxtp_2 _5511_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\ROM_spi_dat_out[1] ),
    .D(_0482_));
 sky130_as_sc_hs__dfxtp_4 _5512_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\ROM_spi_dat_out[2] ),
    .D(_0483_));
 sky130_as_sc_hs__dfxtp_4 _5513_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\ROM_spi_dat_out[3] ),
    .D(_0484_));
 sky130_as_sc_hs__dfxtp_4 _5514_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_14_clk),
    .Q(\ROM_spi_dat_out[4] ),
    .D(_0485_));
 sky130_as_sc_hs__dfxtp_4 _5515_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(\ROM_spi_dat_out[5] ),
    .D(_0486_));
 sky130_as_sc_hs__dfxtp_2 _5516_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(\ROM_spi_dat_out[6] ),
    .D(_0487_));
 sky130_as_sc_hs__dfxtp_2 _5517_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(\ROM_spi_dat_out[7] ),
    .D(_0488_));
 sky130_as_sc_hs__dfxtp_4 _5518_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\ROM_addr_buff[0] ),
    .D(_0489_));
 sky130_as_sc_hs__dfxtp_4 _5519_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\ROM_addr_buff[1] ),
    .D(_0490_));
 sky130_as_sc_hs__dfxtp_4 _5520_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\ROM_addr_buff[2] ),
    .D(_0491_));
 sky130_as_sc_hs__dfxtp_2 _5521_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\ROM_addr_buff[3] ),
    .D(_0492_));
 sky130_as_sc_hs__dfxtp_4 _5522_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\ROM_addr_buff[4] ),
    .D(_0493_));
 sky130_as_sc_hs__dfxtp_2 _5523_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\ROM_addr_buff[5] ),
    .D(_0494_));
 sky130_as_sc_hs__dfxtp_2 _5524_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\ROM_addr_buff[6] ),
    .D(_0495_));
 sky130_as_sc_hs__dfxtp_2 _5525_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\ROM_addr_buff[7] ),
    .D(_0496_));
 sky130_as_sc_hs__dfxtp_2 _5526_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\ROM_addr_buff[8] ),
    .D(_0497_));
 sky130_as_sc_hs__dfxtp_2 _5527_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\ROM_addr_buff[9] ),
    .D(_0498_));
 sky130_as_sc_hs__dfxtp_2 _5528_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\ROM_addr_buff[10] ),
    .D(_0499_));
 sky130_as_sc_hs__dfxtp_2 _5529_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\ROM_addr_buff[11] ),
    .D(_0500_));
 sky130_as_sc_hs__dfxtp_2 _5530_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\last_addr[0] ),
    .D(_0501_));
 sky130_as_sc_hs__dfxtp_2 _5531_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\last_addr[1] ),
    .D(_0502_));
 sky130_as_sc_hs__dfxtp_2 _5532_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\last_addr[2] ),
    .D(_0503_));
 sky130_as_sc_hs__dfxtp_2 _5533_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\last_addr[3] ),
    .D(_0504_));
 sky130_as_sc_hs__dfxtp_2 _5534_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_21_clk),
    .Q(\last_addr[4] ),
    .D(_0505_));
 sky130_as_sc_hs__dfxtp_2 _5535_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\last_addr[5] ),
    .D(_0506_));
 sky130_as_sc_hs__dfxtp_2 _5536_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\last_addr[6] ),
    .D(_0507_));
 sky130_as_sc_hs__dfxtp_2 _5537_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_18_clk),
    .Q(\last_addr[7] ),
    .D(_0508_));
 sky130_as_sc_hs__dfxtp_2 _5538_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\last_addr[8] ),
    .D(_0509_));
 sky130_as_sc_hs__dfxtp_2 _5539_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_19_clk),
    .Q(\last_addr[9] ),
    .D(_0510_));
 sky130_as_sc_hs__dfxtp_2 _5540_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\last_addr[10] ),
    .D(_0511_));
 sky130_as_sc_hs__dfxtp_2 _5541_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_20_clk),
    .Q(\last_addr[11] ),
    .D(_0512_));
 sky130_as_sc_hs__dfxtp_2 _5542_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_13_clk),
    .Q(spi_clkdiv),
    .D(_0513_));
 sky130_as_sc_hs__dfxtp_2 _5543_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_15_clk),
    .Q(\RAM[43][0] ),
    .D(_0514_));
 sky130_as_sc_hs__dfxtp_2 _5544_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_12_clk),
    .Q(\RAM[43][1] ),
    .D(_0515_));
 sky130_as_sc_hs__dfxtp_2 _5545_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_8_clk),
    .Q(\RAM[43][2] ),
    .D(_0516_));
 sky130_as_sc_hs__dfxtp_2 _5546_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[43][3] ),
    .D(_0517_));
 sky130_as_sc_hs__dfxtp_2 _5547_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[43][4] ),
    .D(_0518_));
 sky130_as_sc_hs__dfxtp_2 _5548_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_9_clk),
    .Q(\RAM[43][5] ),
    .D(_0519_));
 sky130_as_sc_hs__dfxtp_2 _5549_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[9][0] ),
    .D(_0520_));
 sky130_as_sc_hs__dfxtp_2 _5550_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_26_clk),
    .Q(\RAM[9][1] ),
    .D(_0521_));
 sky130_as_sc_hs__dfxtp_2 _5551_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[9][2] ),
    .D(_0522_));
 sky130_as_sc_hs__dfxtp_2 _5552_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_31_clk),
    .Q(\RAM[9][3] ),
    .D(_0523_));
 sky130_as_sc_hs__dfxtp_2 _5553_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[9][4] ),
    .D(_0524_));
 sky130_as_sc_hs__dfxtp_2 _5554_ (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .CLK(clknet_leaf_27_clk),
    .Q(\RAM[9][5] ),
    .D(_0525_));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_0_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_0_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__tiel tt_um_sky130_as_sc_hs_164 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ZERO(net164));
 sky130_as_sc_hs__tieh tt_um_sky130_as_sc_hs_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ONE(net165));
 sky130_as_sc_hs__buff_8 _5558_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(CS_ROM),
    .Y(uio_out[7]));
 sky130_as_sc_hs__buff_8 _5559_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ROM_DO),
    .Y(uo_out[6]));
 sky130_as_sc_hs__buff_8 _5560_ (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(SCLK_ROM),
    .Y(uo_out[7]));
 sky130_as_sc_hs__hcf_10 hcf_1 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .HCF(HCF));
 sky130_as_sc_hs__hcf_10 hcf_2 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .HCF(HCF));
 sky130_as_sc_hs__hcf_10 hcf_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .HCF(HCF));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_0_Right_0 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_1_Right_1 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_2_Right_2 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_3_Right_3 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_4_Right_4 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_5_Right_5 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_6_Right_6 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_7_Right_7 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_8_Right_8 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_9_Right_9 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_10_Right_10 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_11_Right_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_12_Right_12 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_13_Right_13 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_14_Right_14 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_15_Right_15 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_16_Right_16 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_17_Right_17 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_18_Right_18 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_19_Right_19 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_20_Right_20 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_21_Right_21 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_22_Right_22 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_23_Right_23 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_24_Right_24 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_25_Right_25 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_26_Right_26 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_27_Right_27 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_28_Right_28 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_29_Right_29 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_30_Right_30 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_31_Right_31 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_32_Right_32 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_33_Right_33 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_34_Right_34 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_35_Right_35 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_36_Right_36 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_37_Right_37 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_38_Right_38 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_39_Right_39 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_40_Right_40 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_41_Right_41 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_42_Right_42 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_43_Right_43 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_44_Right_44 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_45_Right_45 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_46_Right_46 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_47_Right_47 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_48_Right_48 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_49_Right_49 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_50_Right_50 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_51_Right_51 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_52_Right_52 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_53_Right_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_54_Right_54 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_55_Right_55 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_56_Right_56 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_57_Right_57 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_58_Right_58 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_59_Right_59 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_60_Right_60 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_61_Right_61 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_62_Right_62 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_63_Right_63 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_64_Right_64 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_65_Right_65 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_66_Right_66 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_67_Right_67 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_68_Right_68 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_69_Right_69 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_70_Right_70 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_71_Right_71 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_72_Right_72 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_73_Right_73 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_74_Right_74 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_75_Right_75 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_76_Right_76 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_77_Right_77 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_78_Right_78 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_79_Right_79 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_80_Right_80 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_0_Left_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_1_Left_82 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_2_Left_83 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_3_Left_84 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_4_Left_85 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_5_Left_86 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_6_Left_87 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_7_Left_88 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_8_Left_89 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_9_Left_90 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_10_Left_91 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_11_Left_92 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_12_Left_93 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_13_Left_94 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_14_Left_95 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_15_Left_96 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_16_Left_97 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_17_Left_98 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_18_Left_99 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_19_Left_100 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_20_Left_101 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_21_Left_102 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_22_Left_103 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_23_Left_104 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_24_Left_105 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_25_Left_106 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_26_Left_107 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_27_Left_108 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_28_Left_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_29_Left_110 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_30_Left_111 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_31_Left_112 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_32_Left_113 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_33_Left_114 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_34_Left_115 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_35_Left_116 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_36_Left_117 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_37_Left_118 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_38_Left_119 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_39_Left_120 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_40_Left_121 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_41_Left_122 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_42_Left_123 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_43_Left_124 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_44_Left_125 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_45_Left_126 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_46_Left_127 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_47_Left_128 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_48_Left_129 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_49_Left_130 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_50_Left_131 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_51_Left_132 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_52_Left_133 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_53_Left_134 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_54_Left_135 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_55_Left_136 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_56_Left_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_57_Left_138 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_58_Left_139 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_59_Left_140 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_60_Left_141 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_61_Left_142 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_62_Left_143 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_63_Left_144 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_64_Left_145 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_65_Left_146 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_66_Left_147 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_67_Left_148 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_68_Left_149 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_69_Left_150 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_70_Left_151 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_71_Left_152 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_72_Left_153 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_73_Left_154 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_74_Left_155 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_75_Left_156 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_76_Left_157 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_77_Left_158 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_78_Left_159 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_79_Left_160 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 PHY_EDGE_ROW_80_Left_161 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_162 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_163 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_164 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_165 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_166 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_167 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_168 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_169 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_170 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_171 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_172 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_173 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_174 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_175 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_176 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_177 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_178 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_179 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_180 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_181 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_182 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_183 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_184 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_185 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_0_186 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_187 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_188 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_189 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_190 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_191 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_192 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_193 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_194 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_195 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_196 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_197 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_1_198 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_199 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_200 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_201 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_202 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_203 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_204 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_205 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_206 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_207 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_208 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_209 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_210 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_2_211 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_212 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_213 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_214 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_215 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_216 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_217 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_218 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_219 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_220 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_221 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_222 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_3_223 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_224 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_225 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_226 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_227 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_228 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_229 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_230 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_231 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_232 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_233 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_234 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_235 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_4_236 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_237 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_238 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_239 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_240 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_241 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_242 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_243 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_244 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_245 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_246 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_247 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_5_248 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_249 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_250 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_251 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_252 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_253 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_254 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_255 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_256 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_257 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_258 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_259 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_260 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_6_261 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_262 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_263 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_264 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_265 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_266 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_267 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_268 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_269 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_270 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_271 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_272 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_7_273 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_274 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_275 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_276 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_277 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_278 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_279 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_280 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_281 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_282 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_283 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_284 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_285 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_8_286 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_287 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_288 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_289 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_290 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_291 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_292 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_293 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_294 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_295 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_296 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_297 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_9_298 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_299 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_300 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_301 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_302 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_303 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_304 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_305 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_306 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_307 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_308 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_309 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_310 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_10_311 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_312 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_313 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_314 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_315 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_316 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_317 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_318 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_319 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_320 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_321 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_322 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_11_323 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_324 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_325 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_326 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_327 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_328 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_329 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_330 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_331 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_332 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_333 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_334 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_335 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_12_336 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_337 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_338 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_339 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_340 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_341 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_342 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_343 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_344 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_345 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_346 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_347 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_13_348 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_349 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_350 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_351 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_352 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_353 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_354 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_355 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_356 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_357 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_358 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_359 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_360 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_14_361 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_362 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_363 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_364 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_365 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_366 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_367 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_368 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_369 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_370 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_371 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_372 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_15_373 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_374 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_375 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_376 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_377 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_378 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_379 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_380 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_381 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_382 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_383 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_384 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_385 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_16_386 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_387 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_388 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_389 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_390 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_391 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_392 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_393 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_394 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_395 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_396 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_397 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_17_398 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_399 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_400 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_401 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_402 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_403 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_404 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_405 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_406 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_407 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_408 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_409 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_410 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_18_411 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_412 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_413 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_414 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_415 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_416 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_417 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_418 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_419 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_420 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_421 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_422 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_19_423 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_424 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_425 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_426 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_427 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_428 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_429 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_430 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_431 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_432 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_433 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_434 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_435 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_20_436 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_437 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_438 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_439 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_440 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_441 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_442 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_443 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_444 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_445 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_446 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_447 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_21_448 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_449 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_450 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_451 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_452 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_453 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_454 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_455 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_456 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_457 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_458 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_459 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_460 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_22_461 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_462 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_463 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_464 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_465 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_466 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_467 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_468 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_469 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_470 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_471 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_472 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_23_473 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_474 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_475 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_476 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_477 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_478 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_479 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_480 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_481 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_482 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_483 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_484 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_485 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_24_486 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_487 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_488 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_489 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_490 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_491 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_492 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_493 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_494 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_495 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_496 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_497 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_25_498 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_499 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_500 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_501 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_502 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_503 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_504 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_505 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_506 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_507 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_508 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_509 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_510 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_26_511 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_512 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_513 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_514 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_515 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_516 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_517 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_518 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_519 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_520 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_521 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_522 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_27_523 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_524 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_525 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_526 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_527 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_528 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_529 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_530 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_531 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_532 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_533 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_534 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_535 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_28_536 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_537 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_538 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_539 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_540 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_541 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_542 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_543 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_544 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_545 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_546 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_547 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_29_548 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_549 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_550 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_551 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_552 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_553 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_554 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_555 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_556 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_557 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_558 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_559 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_560 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_30_561 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_562 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_563 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_564 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_565 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_566 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_567 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_568 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_569 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_570 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_571 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_572 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_31_573 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_574 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_575 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_576 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_577 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_578 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_579 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_580 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_581 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_582 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_583 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_584 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_585 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_32_586 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_587 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_588 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_589 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_590 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_591 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_592 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_593 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_594 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_595 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_596 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_597 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_33_598 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_599 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_600 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_601 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_602 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_603 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_604 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_605 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_606 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_607 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_608 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_609 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_610 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_34_611 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_612 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_613 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_614 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_615 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_616 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_617 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_618 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_619 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_620 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_621 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_622 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_35_623 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_624 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_625 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_626 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_627 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_628 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_629 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_630 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_631 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_632 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_633 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_634 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_635 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_36_636 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_637 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_638 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_639 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_640 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_641 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_642 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_643 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_644 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_645 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_646 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_647 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_37_648 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_649 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_650 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_651 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_652 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_653 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_654 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_655 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_656 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_657 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_658 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_659 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_660 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_38_661 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_662 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_663 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_664 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_665 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_666 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_667 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_668 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_669 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_670 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_671 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_672 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_39_673 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_674 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_675 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_676 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_677 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_678 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_679 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_680 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_681 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_682 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_683 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_684 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_685 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_40_686 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_687 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_688 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_689 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_690 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_691 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_692 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_693 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_694 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_695 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_696 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_697 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_41_698 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_699 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_700 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_701 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_702 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_703 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_704 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_705 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_706 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_707 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_708 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_709 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_710 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_42_711 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_712 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_713 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_714 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_715 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_716 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_717 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_718 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_719 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_720 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_721 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_722 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_43_723 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_724 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_725 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_726 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_727 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_728 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_729 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_730 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_731 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_732 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_733 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_734 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_735 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_44_736 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_737 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_738 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_739 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_740 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_741 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_742 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_743 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_744 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_745 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_746 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_747 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_45_748 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_749 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_750 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_751 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_752 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_753 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_754 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_755 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_756 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_757 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_758 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_759 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_760 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_46_761 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_762 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_763 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_764 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_765 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_766 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_767 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_768 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_769 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_770 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_771 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_772 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_47_773 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_774 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_775 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_776 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_777 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_778 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_779 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_780 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_781 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_782 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_783 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_784 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_785 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_48_786 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_787 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_788 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_789 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_790 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_791 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_792 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_793 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_794 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_795 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_796 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_797 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_49_798 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_799 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_800 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_801 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_802 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_803 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_804 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_805 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_806 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_807 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_808 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_809 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_810 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_50_811 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_812 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_813 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_814 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_815 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_816 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_817 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_818 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_819 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_820 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_821 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_822 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_51_823 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_824 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_825 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_826 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_827 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_828 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_829 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_830 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_831 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_832 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_833 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_834 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_835 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_52_836 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_837 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_838 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_839 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_840 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_841 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_842 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_843 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_844 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_845 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_846 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_847 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_53_848 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_849 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_850 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_851 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_852 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_853 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_854 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_855 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_856 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_857 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_858 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_859 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_860 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_54_861 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_862 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_863 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_864 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_865 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_866 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_867 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_868 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_869 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_870 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_871 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_872 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_55_873 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_874 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_875 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_876 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_877 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_878 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_879 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_880 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_881 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_882 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_883 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_884 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_885 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_56_886 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_887 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_888 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_889 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_890 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_891 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_892 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_893 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_894 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_895 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_896 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_897 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_57_898 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_899 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_900 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_901 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_902 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_903 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_904 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_905 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_906 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_907 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_908 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_909 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_910 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_58_911 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_912 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_913 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_914 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_915 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_916 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_917 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_918 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_919 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_920 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_921 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_922 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_59_923 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_924 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_925 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_926 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_927 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_928 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_929 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_930 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_931 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_932 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_933 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_934 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_935 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_60_936 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_937 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_938 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_939 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_940 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_941 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_942 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_943 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_944 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_945 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_946 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_947 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_61_948 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_949 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_950 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_951 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_952 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_953 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_954 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_955 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_956 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_957 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_958 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_959 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_960 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_62_961 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_962 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_963 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_964 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_965 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_966 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_967 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_968 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_969 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_970 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_971 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_972 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_63_973 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_974 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_975 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_976 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_977 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_978 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_979 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_980 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_981 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_982 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_983 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_984 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_985 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_64_986 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_987 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_988 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_989 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_990 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_991 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_992 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_993 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_994 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_995 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_996 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_997 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_65_998 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_999 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1000 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1001 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1002 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1003 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1004 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1005 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1006 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1007 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1008 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1009 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1010 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_66_1011 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1012 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1013 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1014 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1015 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1016 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1017 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1018 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1019 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1020 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1021 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1022 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_67_1023 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1024 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1025 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1026 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1027 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1028 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1029 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1030 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1031 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1032 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1033 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1034 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1035 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_68_1036 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1037 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1038 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1039 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1040 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1041 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1042 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1043 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1044 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1045 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1046 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1047 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_69_1048 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1049 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1050 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1051 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1052 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1053 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1054 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1055 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1056 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1057 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1058 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1059 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1060 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_70_1061 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1062 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1063 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1064 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1065 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1066 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1067 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1068 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1069 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1070 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1071 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1072 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_71_1073 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1074 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1075 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1076 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1077 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1078 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1079 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1080 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1081 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1082 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1083 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1084 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1085 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_72_1086 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1087 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1088 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1089 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1090 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1091 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1092 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1093 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1094 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1095 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1096 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1097 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_73_1098 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1099 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1100 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1101 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1102 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1103 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1104 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1105 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1106 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1107 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1108 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1109 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1110 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_74_1111 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1112 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1113 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1114 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1115 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1116 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1117 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1118 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1119 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1120 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1121 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1122 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_75_1123 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1124 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1125 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1126 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1127 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1128 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1129 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1130 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1131 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1132 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1133 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1134 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1135 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_76_1136 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1137 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1138 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1139 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1140 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1141 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1142 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1143 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1144 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1145 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1146 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1147 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_77_1148 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1149 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1150 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1151 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1152 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1153 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1154 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1155 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1156 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1157 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1158 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1159 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1160 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_78_1161 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1162 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1163 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1164 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1165 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1166 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1167 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1168 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1169 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1170 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1171 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1172 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_79_1173 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1174 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1175 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1176 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1177 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1178 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1179 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1180 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1181 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1182 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1183 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1184 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1185 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1186 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1187 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1188 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1189 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1190 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1191 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1192 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1193 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1194 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1195 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1196 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1197 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__tap_1 TAP_TAPCELL_ROW_80_1198 (.VPB(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__buff_2 input1 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(rst_n),
    .Y(net1));
 sky130_as_sc_hs__buff_2 input2 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[0]),
    .Y(net2));
 sky130_as_sc_hs__buff_2 input3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[1]),
    .Y(net3));
 sky130_as_sc_hs__buff_2 input4 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[2]),
    .Y(net4));
 sky130_as_sc_hs__buff_2 input5 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[3]),
    .Y(net5));
 sky130_as_sc_hs__buff_2 input6 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[4]),
    .Y(net6));
 sky130_as_sc_hs__buff_2 input7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[5]),
    .Y(net7));
 sky130_as_sc_hs__buff_2 input8 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[6]),
    .Y(net8));
 sky130_as_sc_hs__buff_2 input9 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(ui_in[7]),
    .Y(net9));
 sky130_as_sc_hs__buff_2 input10 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_in[0]),
    .Y(net10));
 sky130_as_sc_hs__buff_2 input11 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_in[1]),
    .Y(net11));
 sky130_as_sc_hs__buff_2 input12 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_in[2]),
    .Y(net12));
 sky130_as_sc_hs__buff_2 input13 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_in[3]),
    .Y(net13));
 sky130_as_sc_hs__buff_2 input14 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_in[4]),
    .Y(net14));
 sky130_as_sc_hs__buff_2 input15 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_in[5]),
    .Y(net15));
 sky130_as_sc_hs__buff_2 input16 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(uio_in[6]),
    .Y(net16));
 sky130_as_sc_hs__buff_2 max_cap17 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1862_),
    .Y(net17));
 sky130_as_sc_hs__clkbuff_4 max_cap18 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1736_),
    .Y(net18));
 sky130_as_sc_hs__buff_2 max_cap19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net20),
    .Y(net19));
 sky130_as_sc_hs__buff_2 max_cap20 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1569_),
    .Y(net20));
 sky130_as_sc_hs__buff_2 max_cap21 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_1213_),
    .Y(net21));
 sky130_as_sc_hs__buff_2 wire22 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0785_),
    .Y(net22));
 sky130_as_sc_hs__buff_2 max_cap23 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0586_),
    .Y(net23));
 sky130_as_sc_hs__buff_2 max_cap24 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0746_),
    .Y(net24));
 sky130_as_sc_hs__buff_2 max_cap25 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0700_),
    .Y(net25));
 sky130_as_sc_hs__buff_2 max_cap26 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_0698_),
    .Y(net26));
 sky130_as_sc_hs__clkbuff_4 fanout27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\ROM_addr_buff[9] ),
    .Y(net27));
 sky130_as_sc_hs__buff_2 fanout28 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net30),
    .Y(net28));
 sky130_as_sc_hs__buff_2 fanout29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\insin[5] ),
    .Y(net29));
 sky130_as_sc_hs__buff_2 fanout30 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\insin[5] ),
    .Y(net30));
 sky130_as_sc_hs__clkbuff_4 fanout31 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net34),
    .Y(net31));
 sky130_as_sc_hs__clkbuff_4 fanout32 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net33),
    .Y(net32));
 sky130_as_sc_hs__buff_2 fanout33 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net34),
    .Y(net33));
 sky130_as_sc_hs__buff_2 fanout34 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\insin[4] ),
    .Y(net34));
 sky130_as_sc_hs__clkbuff_4 fanout35 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\insin[3] ),
    .Y(net35));
 sky130_as_sc_hs__buff_2 fanout36 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\insin[3] ),
    .Y(net36));
 sky130_as_sc_hs__buff_4 fanout37 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net38),
    .Y(net37));
 sky130_as_sc_hs__buff_2 fanout38 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net39),
    .Y(net38));
 sky130_as_sc_hs__buff_4 fanout39 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\insin[2] ),
    .Y(net39));
 sky130_as_sc_hs__clkbuff_4 fanout40 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net44),
    .Y(net40));
 sky130_as_sc_hs__clkbuff_4 fanout41 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net42),
    .Y(net41));
 sky130_as_sc_hs__buff_2 fanout42 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net43),
    .Y(net42));
 sky130_as_sc_hs__clkbuff_4 fanout43 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net44),
    .Y(net43));
 sky130_as_sc_hs__buff_2 fanout44 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\insin[1] ),
    .Y(net44));
 sky130_as_sc_hs__buff_4 fanout45 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net47),
    .Y(net45));
 sky130_as_sc_hs__buff_2 fanout46 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net47),
    .Y(net46));
 sky130_as_sc_hs__clkbuff_4 fanout47 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\insin[0] ),
    .Y(net47));
 sky130_as_sc_hs__buff_8 fanout48 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\insin[0] ),
    .Y(net48));
 sky130_as_sc_hs__clkbuff_4 fanout49 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net50),
    .Y(net49));
 sky130_as_sc_hs__buff_2 fanout50 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[4] ),
    .Y(net50));
 sky130_as_sc_hs__buff_4 fanout51 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[4] ),
    .Y(net51));
 sky130_as_sc_hs__clkbuff_4 fanout52 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net53),
    .Y(net52));
 sky130_as_sc_hs__buff_2 fanout53 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net54),
    .Y(net53));
 sky130_as_sc_hs__buff_4 fanout54 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net55),
    .Y(net54));
 sky130_as_sc_hs__clkbuff_4 fanout55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[3] ),
    .Y(net55));
 sky130_as_sc_hs__buff_4 fanout56 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net57),
    .Y(net56));
 sky130_as_sc_hs__buff_2 fanout57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net63),
    .Y(net57));
 sky130_as_sc_hs__clkbuff_4 fanout58 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net60),
    .Y(net58));
 sky130_as_sc_hs__buff_2 fanout59 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net60),
    .Y(net59));
 sky130_as_sc_hs__buff_4 fanout60 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net63),
    .Y(net60));
 sky130_as_sc_hs__buff_4 fanout61 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net63),
    .Y(net61));
 sky130_as_sc_hs__buff_8 fanout62 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net63),
    .Y(net62));
 sky130_as_sc_hs__clkbuff_4 fanout63 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[2] ),
    .Y(net63));
 sky130_as_sc_hs__buff_4 fanout64 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net66),
    .Y(net64));
 sky130_as_sc_hs__buff_2 fanout65 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net66),
    .Y(net65));
 sky130_as_sc_hs__buff_4 fanout66 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net69),
    .Y(net66));
 sky130_as_sc_hs__buff_4 fanout67 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net68),
    .Y(net67));
 sky130_as_sc_hs__buff_4 fanout68 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net69),
    .Y(net68));
 sky130_as_sc_hs__buff_2 fanout69 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net74),
    .Y(net69));
 sky130_as_sc_hs__buff_4 fanout70 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net71),
    .Y(net70));
 sky130_as_sc_hs__buff_4 fanout71 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net72),
    .Y(net71));
 sky130_as_sc_hs__buff_4 fanout72 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net74),
    .Y(net72));
 sky130_as_sc_hs__buff_2 fanout73 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net74),
    .Y(net73));
 sky130_as_sc_hs__buff_2 fanout74 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net89),
    .Y(net74));
 sky130_as_sc_hs__buff_4 fanout75 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net77),
    .Y(net75));
 sky130_as_sc_hs__buff_2 fanout76 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net77),
    .Y(net76));
 sky130_as_sc_hs__buff_4 fanout77 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net83),
    .Y(net77));
 sky130_as_sc_hs__buff_4 fanout78 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net82),
    .Y(net78));
 sky130_as_sc_hs__buff_2 fanout79 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net82),
    .Y(net79));
 sky130_as_sc_hs__buff_4 fanout80 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net82),
    .Y(net80));
 sky130_as_sc_hs__buff_2 fanout81 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net82),
    .Y(net81));
 sky130_as_sc_hs__buff_2 fanout82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net83),
    .Y(net82));
 sky130_as_sc_hs__buff_2 fanout83 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net89),
    .Y(net83));
 sky130_as_sc_hs__buff_4 fanout84 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net85),
    .Y(net84));
 sky130_as_sc_hs__buff_4 fanout85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net88),
    .Y(net85));
 sky130_as_sc_hs__buff_4 fanout86 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net87),
    .Y(net86));
 sky130_as_sc_hs__buff_4 fanout87 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net88),
    .Y(net87));
 sky130_as_sc_hs__buff_2 fanout88 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net89),
    .Y(net88));
 sky130_as_sc_hs__buff_2 fanout89 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[1] ),
    .Y(net89));
 sky130_as_sc_hs__buff_4 fanout90 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net95),
    .Y(net90));
 sky130_as_sc_hs__buff_2 fanout91 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net95),
    .Y(net91));
 sky130_as_sc_hs__buff_4 fanout92 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net95),
    .Y(net92));
 sky130_as_sc_hs__buff_4 fanout93 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net95),
    .Y(net93));
 sky130_as_sc_hs__clkbuff_4 fanout94 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net95),
    .Y(net94));
 sky130_as_sc_hs__buff_2 fanout95 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net103),
    .Y(net95));
 sky130_as_sc_hs__buff_4 fanout96 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net100),
    .Y(net96));
 sky130_as_sc_hs__buff_4 fanout97 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net100),
    .Y(net97));
 sky130_as_sc_hs__buff_4 fanout98 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net99),
    .Y(net98));
 sky130_as_sc_hs__buff_4 fanout99 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net100),
    .Y(net99));
 sky130_as_sc_hs__buff_2 fanout100 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net103),
    .Y(net100));
 sky130_as_sc_hs__buff_4 fanout101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net103),
    .Y(net101));
 sky130_as_sc_hs__buff_2 fanout102 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net103),
    .Y(net102));
 sky130_as_sc_hs__buff_2 fanout103 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[1] ),
    .Y(net103));
 sky130_as_sc_hs__buff_4 fanout104 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net108),
    .Y(net104));
 sky130_as_sc_hs__clkbuff_4 fanout105 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net108),
    .Y(net105));
 sky130_as_sc_hs__buff_4 fanout106 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net108),
    .Y(net106));
 sky130_as_sc_hs__buff_2 fanout107 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net108),
    .Y(net107));
 sky130_as_sc_hs__buff_2 fanout108 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net118),
    .Y(net108));
 sky130_as_sc_hs__buff_4 fanout109 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net111),
    .Y(net109));
 sky130_as_sc_hs__buff_4 fanout110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net111),
    .Y(net110));
 sky130_as_sc_hs__clkbuff_4 fanout111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net118),
    .Y(net111));
 sky130_as_sc_hs__buff_4 fanout112 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net113),
    .Y(net112));
 sky130_as_sc_hs__buff_8 fanout113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net117),
    .Y(net113));
 sky130_as_sc_hs__buff_4 fanout114 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net115),
    .Y(net114));
 sky130_as_sc_hs__clkbuff_4 fanout115 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net116),
    .Y(net115));
 sky130_as_sc_hs__buff_2 fanout116 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net117),
    .Y(net116));
 sky130_as_sc_hs__clkbuff_4 fanout117 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net118),
    .Y(net117));
 sky130_as_sc_hs__buff_2 fanout118 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[0] ),
    .Y(net118));
 sky130_as_sc_hs__buff_4 fanout119 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net121),
    .Y(net119));
 sky130_as_sc_hs__buff_8 fanout120 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net121),
    .Y(net120));
 sky130_as_sc_hs__clkbuff_4 fanout121 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net123),
    .Y(net121));
 sky130_as_sc_hs__clkbuff_4 fanout122 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net123),
    .Y(net122));
 sky130_as_sc_hs__buff_2 fanout123 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[0] ),
    .Y(net123));
 sky130_as_sc_hs__clkbuff_4 fanout124 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\A[5] ),
    .Y(net124));
 sky130_as_sc_hs__buff_2 fanout125 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\A[5] ),
    .Y(net125));
 sky130_as_sc_hs__clkbuff_4 fanout126 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\A[4] ),
    .Y(net126));
 sky130_as_sc_hs__clkbuff_4 fanout127 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\A[4] ),
    .Y(net127));
 sky130_as_sc_hs__clkbuff_4 fanout128 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net129),
    .Y(net128));
 sky130_as_sc_hs__clkbuff_4 fanout129 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\A[2] ),
    .Y(net129));
 sky130_as_sc_hs__clkbuff_4 fanout130 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net131),
    .Y(net130));
 sky130_as_sc_hs__buff_2 fanout131 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\A[1] ),
    .Y(net131));
 sky130_as_sc_hs__clkbuff_4 fanout132 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\A[0] ),
    .Y(net132));
 sky130_as_sc_hs__buff_2 fanout133 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\A[0] ),
    .Y(net133));
 sky130_as_sc_hs__buff_4 fanout134 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net137),
    .Y(net134));
 sky130_as_sc_hs__clkbuff_4 fanout135 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net136),
    .Y(net135));
 sky130_as_sc_hs__clkbuff_4 fanout136 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net137),
    .Y(net136));
 sky130_as_sc_hs__buff_2 fanout137 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\instr_cycle[2] ),
    .Y(net137));
 sky130_as_sc_hs__clkbuff_4 fanout138 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\instr_cycle[0] ),
    .Y(net138));
 sky130_as_sc_hs__buff_2 fanout139 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\instr_cycle[0] ),
    .Y(net139));
 sky130_as_sc_hs__buff_4 fanout140 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net142),
    .Y(net140));
 sky130_as_sc_hs__buff_4 fanout141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[5] ),
    .Y(net141));
 sky130_as_sc_hs__buff_2 fanout142 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\MAR[5] ),
    .Y(net142));
 sky130_as_sc_hs__clkbuff_4 fanout143 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\mem_cycle[2] ),
    .Y(net143));
 sky130_as_sc_hs__clkbuff_4 fanout144 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net145),
    .Y(net144));
 sky130_as_sc_hs__clkbuff_4 fanout145 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\mem_cycle[0] ),
    .Y(net145));
 sky130_as_sc_hs__buff_2 fanout146 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net147),
    .Y(net146));
 sky130_as_sc_hs__buff_2 fanout147 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net148),
    .Y(net147));
 sky130_as_sc_hs__buff_2 fanout148 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net162),
    .Y(net148));
 sky130_as_sc_hs__buff_2 fanout149 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net153),
    .Y(net149));
 sky130_as_sc_hs__buff_2 fanout150 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net153),
    .Y(net150));
 sky130_as_sc_hs__buff_2 fanout151 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net152),
    .Y(net151));
 sky130_as_sc_hs__buff_2 fanout152 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net153),
    .Y(net152));
 sky130_as_sc_hs__buff_2 fanout153 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net162),
    .Y(net153));
 sky130_as_sc_hs__buff_2 fanout154 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net156),
    .Y(net154));
 sky130_as_sc_hs__buff_2 fanout155 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net156),
    .Y(net155));
 sky130_as_sc_hs__buff_2 fanout156 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net161),
    .Y(net156));
 sky130_as_sc_hs__clkbuff_4 fanout157 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net161),
    .Y(net157));
 sky130_as_sc_hs__buff_2 fanout158 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net160),
    .Y(net158));
 sky130_as_sc_hs__buff_2 fanout159 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net160),
    .Y(net159));
 sky130_as_sc_hs__buff_4 fanout160 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net161),
    .Y(net160));
 sky130_as_sc_hs__buff_2 fanout161 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net162),
    .Y(net161));
 sky130_as_sc_hs__buff_2 fanout162 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(net1),
    .Y(net162));
 sky130_as_sc_hs__tiel tt_um_sky130_as_sc_hs_163 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .ZERO(net163));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_1_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_1_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_2_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_2_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_3_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_3_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_4_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_4_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_5_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_5_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_6_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_6_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_7_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_7_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_8_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_8_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_9_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_9_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_10_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_10_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_11_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_11_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_12_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_12_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_13_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_13_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_14_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_14_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_15_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_15_clk),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_16_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_16_clk),
    .A(clknet_2_2__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_17_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_17_clk),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_18_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_18_clk),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_19_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_19_clk),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_20_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_20_clk),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_21_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_21_clk),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_22_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_22_clk),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_23_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_23_clk),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_24_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_24_clk),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_25_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_25_clk),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_26_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_26_clk),
    .A(clknet_2_2__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_27_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_27_clk),
    .A(clknet_2_2__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_28_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_28_clk),
    .A(clknet_2_2__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_29_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_29_clk),
    .A(clknet_2_2__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_30_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_30_clk),
    .A(clknet_2_2__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_31_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_31_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_32_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_32_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_33_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_33_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_34_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_34_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_35_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_35_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_8 clkbuf_leaf_36_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .Y(clknet_leaf_36_clk),
    .A(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_11 clkbuf_0_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clk),
    .Y(clknet_0_clk));
 sky130_as_sc_hs__clkbuff_11 clkbuf_2_0__f_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_0_clk),
    .Y(clknet_2_0__leaf_clk));
 sky130_as_sc_hs__clkbuff_11 clkbuf_2_1__f_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_0_clk),
    .Y(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__clkbuff_11 clkbuf_2_2__f_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_0_clk),
    .Y(clknet_2_2__leaf_clk));
 sky130_as_sc_hs__clkbuff_11 clkbuf_2_3__f_clk (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_0_clk),
    .Y(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__inv_4 clkload0 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_2_1__leaf_clk));
 sky130_as_sc_hs__inv_6 clkload1 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_2_2__leaf_clk));
 sky130_as_sc_hs__inv_6 clkload2 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_2_3__leaf_clk));
 sky130_as_sc_hs__clkbuff_4 clkload3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_leaf_0_clk));
 sky130_as_sc_hs__inv_6 clkload4 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_1_clk));
 sky130_as_sc_hs__inv_4 clkload5 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_2_clk));
 sky130_as_sc_hs__inv_4 clkload6 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_3_clk));
 sky130_as_sc_hs__clkbuff_4 clkload7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_leaf_4_clk));
 sky130_as_sc_hs__inv_6 clkload8 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_5_clk));
 sky130_as_sc_hs__clkbuff_4 clkload9 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_leaf_31_clk));
 sky130_as_sc_hs__inv_6 clkload10 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_32_clk));
 sky130_as_sc_hs__inv_6 clkload11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_33_clk));
 sky130_as_sc_hs__inv_4 clkload12 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_35_clk));
 sky130_as_sc_hs__inv_6 clkload13 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_36_clk));
 sky130_as_sc_hs__inv_2 clkload14 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_6_clk));
 sky130_as_sc_hs__clkbuff_4 clkload15 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_leaf_7_clk));
 sky130_as_sc_hs__inv_4 clkload16 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_8_clk));
 sky130_as_sc_hs__inv_2 clkload17 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_9_clk));
 sky130_as_sc_hs__clkbuff_4 clkload18 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_leaf_10_clk));
 sky130_as_sc_hs__clkbuff_4 clkload19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(clknet_leaf_11_clk));
 sky130_as_sc_hs__inv_4 clkload20 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_13_clk));
 sky130_as_sc_hs__inv_4 clkload21 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_14_clk));
 sky130_as_sc_hs__inv_6 clkload22 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_15_clk));
 sky130_as_sc_hs__inv_4 clkload23 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_16_clk));
 sky130_as_sc_hs__inv_4 clkload24 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_26_clk));
 sky130_as_sc_hs__inv_6 clkload25 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_27_clk));
 sky130_as_sc_hs__inv_6 clkload26 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_28_clk));
 sky130_as_sc_hs__inv_6 clkload27 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_29_clk));
 sky130_as_sc_hs__inv_6 clkload28 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_17_clk));
 sky130_as_sc_hs__inv_4 clkload29 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_18_clk));
 sky130_as_sc_hs__inv_6 clkload30 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_20_clk));
 sky130_as_sc_hs__inv_4 clkload31 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_21_clk));
 sky130_as_sc_hs__inv_2 clkload32 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_22_clk));
 sky130_as_sc_hs__inv_6 clkload33 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_23_clk));
 sky130_as_sc_hs__inv_6 clkload34 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_24_clk));
 sky130_as_sc_hs__inv_6 clkload35 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR),
    .A(clknet_leaf_25_clk));
 sky130_as_sc_hs__buff_2 hold1 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\B[2] ),
    .Y(net166));
 sky130_as_sc_hs__buff_2 hold2 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2138_),
    .Y(net167));
 sky130_as_sc_hs__buff_2 hold3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\ROM_dest[0] ),
    .Y(net168));
 sky130_as_sc_hs__buff_2 hold4 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\B[3] ),
    .Y(net169));
 sky130_as_sc_hs__buff_2 hold5 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(spi_clkdiv),
    .Y(net170));
 sky130_as_sc_hs__buff_2 hold6 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2499_),
    .Y(net171));
 sky130_as_sc_hs__buff_2 hold7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(needs_irupt),
    .Y(net172));
 sky130_as_sc_hs__buff_2 hold8 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2358_),
    .Y(net173));
 sky130_as_sc_hs__buff_2 hold9 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_MAR[3] ),
    .Y(net174));
 sky130_as_sc_hs__buff_2 hold10 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\imm_buff[2] ),
    .Y(net175));
 sky130_as_sc_hs__buff_2 hold11 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[10] ),
    .Y(net176));
 sky130_as_sc_hs__buff_2 hold12 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_P[3] ),
    .Y(net177));
 sky130_as_sc_hs__buff_2 hold13 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[11] ),
    .Y(net178));
 sky130_as_sc_hs__buff_2 hold14 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[43][0] ),
    .Y(net179));
 sky130_as_sc_hs__buff_2 hold15 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_P[0] ),
    .Y(net180));
 sky130_as_sc_hs__buff_2 hold16 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[9] ),
    .Y(net181));
 sky130_as_sc_hs__buff_2 hold17 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\PC[2] ),
    .Y(net182));
 sky130_as_sc_hs__buff_2 hold18 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[8] ),
    .Y(net183));
 sky130_as_sc_hs__buff_2 hold19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\imm_buff[1] ),
    .Y(net184));
 sky130_as_sc_hs__buff_2 hold20 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[7] ),
    .Y(net185));
 sky130_as_sc_hs__buff_2 hold21 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[6] ),
    .Y(net186));
 sky130_as_sc_hs__buff_2 hold22 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2321_),
    .Y(net187));
 sky130_as_sc_hs__buff_2 hold23 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[22][3] ),
    .Y(net188));
 sky130_as_sc_hs__buff_2 hold24 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_MAR[2] ),
    .Y(net189));
 sky130_as_sc_hs__buff_2 hold25 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_P[2] ),
    .Y(net190));
 sky130_as_sc_hs__buff_2 hold26 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[43][1] ),
    .Y(net191));
 sky130_as_sc_hs__buff_2 hold27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[57][0] ),
    .Y(net192));
 sky130_as_sc_hs__buff_2 hold28 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[43][2] ),
    .Y(net193));
 sky130_as_sc_hs__buff_2 hold29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_P[5] ),
    .Y(net194));
 sky130_as_sc_hs__buff_2 hold30 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[57][4] ),
    .Y(net195));
 sky130_as_sc_hs__buff_2 hold31 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[16][0] ),
    .Y(net196));
 sky130_as_sc_hs__buff_2 hold32 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[32][2] ),
    .Y(net197));
 sky130_as_sc_hs__buff_2 hold33 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[49][0] ),
    .Y(net198));
 sky130_as_sc_hs__buff_2 hold34 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[56][3] ),
    .Y(net199));
 sky130_as_sc_hs__buff_2 hold35 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[23][0] ),
    .Y(net200));
 sky130_as_sc_hs__buff_2 hold36 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_P[4] ),
    .Y(net201));
 sky130_as_sc_hs__buff_2 hold37 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[25][5] ),
    .Y(net202));
 sky130_as_sc_hs__buff_2 hold38 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[57][5] ),
    .Y(net203));
 sky130_as_sc_hs__buff_2 hold39 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[56][1] ),
    .Y(net204));
 sky130_as_sc_hs__buff_2 hold40 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[2] ),
    .Y(net205));
 sky130_as_sc_hs__buff_2 hold41 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_B[2] ),
    .Y(net206));
 sky130_as_sc_hs__buff_2 hold42 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[34][0] ),
    .Y(net207));
 sky130_as_sc_hs__buff_2 hold43 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[20][0] ),
    .Y(net208));
 sky130_as_sc_hs__buff_2 hold44 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[10][0] ),
    .Y(net209));
 sky130_as_sc_hs__buff_2 hold45 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[14][3] ),
    .Y(net210));
 sky130_as_sc_hs__buff_2 hold46 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[18][0] ),
    .Y(net211));
 sky130_as_sc_hs__buff_2 hold47 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_B[5] ),
    .Y(net212));
 sky130_as_sc_hs__buff_2 hold48 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2343_),
    .Y(net213));
 sky130_as_sc_hs__buff_2 hold49 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[22][1] ),
    .Y(net214));
 sky130_as_sc_hs__buff_2 hold50 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[45][3] ),
    .Y(net215));
 sky130_as_sc_hs__buff_2 hold51 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[31][1] ),
    .Y(net216));
 sky130_as_sc_hs__buff_2 hold52 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[0][1] ),
    .Y(net217));
 sky130_as_sc_hs__buff_2 hold53 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[30][2] ),
    .Y(net218));
 sky130_as_sc_hs__buff_2 hold54 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_B[3] ),
    .Y(net219));
 sky130_as_sc_hs__buff_2 hold55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_A[1] ),
    .Y(net220));
 sky130_as_sc_hs__buff_2 hold56 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[5] ),
    .Y(net221));
 sky130_as_sc_hs__buff_2 hold57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[13][2] ),
    .Y(net222));
 sky130_as_sc_hs__buff_2 hold58 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[36][5] ),
    .Y(net223));
 sky130_as_sc_hs__buff_2 hold59 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[54][3] ),
    .Y(net224));
 sky130_as_sc_hs__buff_2 hold60 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[36][0] ),
    .Y(net225));
 sky130_as_sc_hs__buff_2 hold61 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[33][1] ),
    .Y(net226));
 sky130_as_sc_hs__buff_2 hold62 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[4][0] ),
    .Y(net227));
 sky130_as_sc_hs__buff_2 hold63 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[27][0] ),
    .Y(net228));
 sky130_as_sc_hs__buff_2 hold64 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[62][0] ),
    .Y(net229));
 sky130_as_sc_hs__buff_2 hold65 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[30][0] ),
    .Y(net230));
 sky130_as_sc_hs__buff_2 hold66 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[27][4] ),
    .Y(net231));
 sky130_as_sc_hs__buff_2 hold67 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[31][0] ),
    .Y(net232));
 sky130_as_sc_hs__buff_2 hold68 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[3][2] ),
    .Y(net233));
 sky130_as_sc_hs__buff_2 hold69 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[20][3] ),
    .Y(net234));
 sky130_as_sc_hs__buff_2 hold70 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[42][5] ),
    .Y(net235));
 sky130_as_sc_hs__buff_2 hold71 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[28][1] ),
    .Y(net236));
 sky130_as_sc_hs__buff_2 hold72 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[3][5] ),
    .Y(net237));
 sky130_as_sc_hs__buff_2 hold73 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[12][3] ),
    .Y(net238));
 sky130_as_sc_hs__buff_2 hold74 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[21][3] ),
    .Y(net239));
 sky130_as_sc_hs__buff_2 hold75 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[7][5] ),
    .Y(net240));
 sky130_as_sc_hs__buff_2 hold76 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[48][0] ),
    .Y(net241));
 sky130_as_sc_hs__buff_2 hold77 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[38][5] ),
    .Y(net242));
 sky130_as_sc_hs__buff_2 hold78 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[40][4] ),
    .Y(net243));
 sky130_as_sc_hs__buff_2 hold79 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[61][3] ),
    .Y(net244));
 sky130_as_sc_hs__buff_2 hold80 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_MAR[5] ),
    .Y(net245));
 sky130_as_sc_hs__buff_2 hold81 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[39][0] ),
    .Y(net246));
 sky130_as_sc_hs__buff_2 hold82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[33][2] ),
    .Y(net247));
 sky130_as_sc_hs__buff_2 hold83 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[34][3] ),
    .Y(net248));
 sky130_as_sc_hs__buff_2 hold84 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[11][4] ),
    .Y(net249));
 sky130_as_sc_hs__buff_2 hold85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[61][1] ),
    .Y(net250));
 sky130_as_sc_hs__buff_2 hold86 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[18][1] ),
    .Y(net251));
 sky130_as_sc_hs__buff_2 hold87 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[32][3] ),
    .Y(net252));
 sky130_as_sc_hs__buff_2 hold88 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[24][0] ),
    .Y(net253));
 sky130_as_sc_hs__buff_2 hold89 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[14][0] ),
    .Y(net254));
 sky130_as_sc_hs__buff_2 hold90 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[40][0] ),
    .Y(net255));
 sky130_as_sc_hs__buff_2 hold91 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\imm_buff[0] ),
    .Y(net256));
 sky130_as_sc_hs__buff_2 hold92 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[54][1] ),
    .Y(net257));
 sky130_as_sc_hs__buff_2 hold93 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[10][2] ),
    .Y(net258));
 sky130_as_sc_hs__buff_2 hold94 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[57][1] ),
    .Y(net259));
 sky130_as_sc_hs__buff_2 hold95 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[35][1] ),
    .Y(net260));
 sky130_as_sc_hs__buff_2 hold96 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[51][3] ),
    .Y(net261));
 sky130_as_sc_hs__buff_2 hold97 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[33][5] ),
    .Y(net262));
 sky130_as_sc_hs__buff_2 hold98 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[30][1] ),
    .Y(net263));
 sky130_as_sc_hs__buff_2 hold99 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[26][0] ),
    .Y(net264));
 sky130_as_sc_hs__buff_2 hold100 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[6][3] ),
    .Y(net265));
 sky130_as_sc_hs__buff_2 hold101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[15][2] ),
    .Y(net266));
 sky130_as_sc_hs__buff_2 hold102 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[12][1] ),
    .Y(net267));
 sky130_as_sc_hs__buff_2 hold103 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[26][3] ),
    .Y(net268));
 sky130_as_sc_hs__buff_2 hold104 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[54][2] ),
    .Y(net269));
 sky130_as_sc_hs__buff_2 hold105 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[5][2] ),
    .Y(net270));
 sky130_as_sc_hs__buff_2 hold106 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[25][1] ),
    .Y(net271));
 sky130_as_sc_hs__buff_2 hold107 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[12][4] ),
    .Y(net272));
 sky130_as_sc_hs__buff_2 hold108 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[16][1] ),
    .Y(net273));
 sky130_as_sc_hs__buff_2 hold109 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[15][3] ),
    .Y(net274));
 sky130_as_sc_hs__buff_2 hold110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[9][4] ),
    .Y(net275));
 sky130_as_sc_hs__buff_2 hold111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[6][1] ),
    .Y(net276));
 sky130_as_sc_hs__buff_2 hold112 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[46][1] ),
    .Y(net277));
 sky130_as_sc_hs__buff_2 hold113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[3][4] ),
    .Y(net278));
 sky130_as_sc_hs__buff_2 hold114 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[11][3] ),
    .Y(net279));
 sky130_as_sc_hs__buff_2 hold115 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[11][0] ),
    .Y(net280));
 sky130_as_sc_hs__buff_2 hold116 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[40][3] ),
    .Y(net281));
 sky130_as_sc_hs__buff_2 hold117 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[30][4] ),
    .Y(net282));
 sky130_as_sc_hs__buff_2 hold118 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[44][1] ),
    .Y(net283));
 sky130_as_sc_hs__buff_2 hold119 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[27][1] ),
    .Y(net284));
 sky130_as_sc_hs__buff_2 hold120 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[37][5] ),
    .Y(net285));
 sky130_as_sc_hs__buff_2 hold121 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_A[2] ),
    .Y(net286));
 sky130_as_sc_hs__buff_2 hold122 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[48][2] ),
    .Y(net287));
 sky130_as_sc_hs__buff_2 hold123 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[41][5] ),
    .Y(net288));
 sky130_as_sc_hs__buff_2 hold124 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[33][4] ),
    .Y(net289));
 sky130_as_sc_hs__buff_2 hold125 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[4][5] ),
    .Y(net290));
 sky130_as_sc_hs__buff_2 hold126 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[35][0] ),
    .Y(net291));
 sky130_as_sc_hs__buff_2 hold127 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[15][4] ),
    .Y(net292));
 sky130_as_sc_hs__buff_2 hold128 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[45][0] ),
    .Y(net293));
 sky130_as_sc_hs__buff_2 hold129 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[19][1] ),
    .Y(net294));
 sky130_as_sc_hs__buff_2 hold130 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[52][0] ),
    .Y(net295));
 sky130_as_sc_hs__buff_2 hold131 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[39][5] ),
    .Y(net296));
 sky130_as_sc_hs__buff_2 hold132 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[17][2] ),
    .Y(net297));
 sky130_as_sc_hs__buff_2 hold133 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[42][4] ),
    .Y(net298));
 sky130_as_sc_hs__buff_2 hold134 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[31][3] ),
    .Y(net299));
 sky130_as_sc_hs__buff_2 hold135 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[55][0] ),
    .Y(net300));
 sky130_as_sc_hs__buff_2 hold136 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[28][2] ),
    .Y(net301));
 sky130_as_sc_hs__buff_2 hold137 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[37][1] ),
    .Y(net302));
 sky130_as_sc_hs__buff_2 hold138 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[36][1] ),
    .Y(net303));
 sky130_as_sc_hs__buff_2 hold139 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[44][0] ),
    .Y(net304));
 sky130_as_sc_hs__buff_2 hold140 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[15][0] ),
    .Y(net305));
 sky130_as_sc_hs__buff_2 hold141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[31][4] ),
    .Y(net306));
 sky130_as_sc_hs__buff_2 hold142 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[53][0] ),
    .Y(net307));
 sky130_as_sc_hs__buff_2 hold143 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[21][4] ),
    .Y(net308));
 sky130_as_sc_hs__buff_2 hold144 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[37][2] ),
    .Y(net309));
 sky130_as_sc_hs__buff_2 hold145 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[25][0] ),
    .Y(net310));
 sky130_as_sc_hs__buff_2 hold146 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[48][1] ),
    .Y(net311));
 sky130_as_sc_hs__buff_2 hold147 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[40][5] ),
    .Y(net312));
 sky130_as_sc_hs__buff_2 hold148 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[35][2] ),
    .Y(net313));
 sky130_as_sc_hs__buff_2 hold149 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[41][4] ),
    .Y(net314));
 sky130_as_sc_hs__buff_2 hold150 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[12][5] ),
    .Y(net315));
 sky130_as_sc_hs__buff_2 hold151 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[40][1] ),
    .Y(net316));
 sky130_as_sc_hs__buff_2 hold152 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[19][3] ),
    .Y(net317));
 sky130_as_sc_hs__buff_2 hold153 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[17][0] ),
    .Y(net318));
 sky130_as_sc_hs__buff_2 hold154 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[33][0] ),
    .Y(net319));
 sky130_as_sc_hs__buff_2 hold155 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[27][2] ),
    .Y(net320));
 sky130_as_sc_hs__buff_2 hold156 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[37][4] ),
    .Y(net321));
 sky130_as_sc_hs__buff_2 hold157 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[44][2] ),
    .Y(net322));
 sky130_as_sc_hs__buff_2 hold158 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[37][0] ),
    .Y(net323));
 sky130_as_sc_hs__buff_2 hold159 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[11][2] ),
    .Y(net324));
 sky130_as_sc_hs__buff_2 hold160 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[47][2] ),
    .Y(net325));
 sky130_as_sc_hs__buff_2 hold161 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[49][2] ),
    .Y(net326));
 sky130_as_sc_hs__buff_2 hold162 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[52][4] ),
    .Y(net327));
 sky130_as_sc_hs__buff_2 hold163 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[54][0] ),
    .Y(net328));
 sky130_as_sc_hs__buff_2 hold164 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[53][3] ),
    .Y(net329));
 sky130_as_sc_hs__buff_2 hold165 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[17][3] ),
    .Y(net330));
 sky130_as_sc_hs__buff_2 hold166 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[2][0] ),
    .Y(net331));
 sky130_as_sc_hs__buff_2 hold167 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[46][2] ),
    .Y(net332));
 sky130_as_sc_hs__buff_2 hold168 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_MAR[4] ),
    .Y(net333));
 sky130_as_sc_hs__buff_2 hold169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[23][5] ),
    .Y(net334));
 sky130_as_sc_hs__buff_2 hold170 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[40][2] ),
    .Y(net335));
 sky130_as_sc_hs__buff_2 hold171 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[38][2] ),
    .Y(net336));
 sky130_as_sc_hs__buff_2 hold172 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[21][0] ),
    .Y(net337));
 sky130_as_sc_hs__buff_2 hold173 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[4][3] ),
    .Y(net338));
 sky130_as_sc_hs__buff_2 hold174 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[28][0] ),
    .Y(net339));
 sky130_as_sc_hs__buff_2 hold175 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[20][4] ),
    .Y(net340));
 sky130_as_sc_hs__buff_2 hold176 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[1][4] ),
    .Y(net341));
 sky130_as_sc_hs__buff_2 hold177 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[7][2] ),
    .Y(net342));
 sky130_as_sc_hs__buff_2 hold178 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[24][3] ),
    .Y(net343));
 sky130_as_sc_hs__buff_2 hold179 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[4][1] ),
    .Y(net344));
 sky130_as_sc_hs__buff_2 hold180 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[9][2] ),
    .Y(net345));
 sky130_as_sc_hs__buff_2 hold181 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[26][5] ),
    .Y(net346));
 sky130_as_sc_hs__buff_2 hold182 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[13][4] ),
    .Y(net347));
 sky130_as_sc_hs__buff_2 hold183 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[20][5] ),
    .Y(net348));
 sky130_as_sc_hs__buff_2 hold184 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[6][0] ),
    .Y(net349));
 sky130_as_sc_hs__buff_2 hold185 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[52][2] ),
    .Y(net350));
 sky130_as_sc_hs__buff_2 hold186 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[39][1] ),
    .Y(net351));
 sky130_as_sc_hs__buff_2 hold187 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[45][1] ),
    .Y(net352));
 sky130_as_sc_hs__buff_2 hold188 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[39][4] ),
    .Y(net353));
 sky130_as_sc_hs__buff_2 hold189 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[46][4] ),
    .Y(net354));
 sky130_as_sc_hs__buff_2 hold190 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[44][3] ),
    .Y(net355));
 sky130_as_sc_hs__buff_2 hold191 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[55][1] ),
    .Y(net356));
 sky130_as_sc_hs__buff_2 hold192 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[53][1] ),
    .Y(net357));
 sky130_as_sc_hs__buff_2 hold193 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[57][3] ),
    .Y(net358));
 sky130_as_sc_hs__buff_2 hold194 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[15][5] ),
    .Y(net359));
 sky130_as_sc_hs__buff_2 hold195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[14][5] ),
    .Y(net360));
 sky130_as_sc_hs__buff_2 hold196 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[35][4] ),
    .Y(net361));
 sky130_as_sc_hs__buff_2 hold197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[47][0] ),
    .Y(net362));
 sky130_as_sc_hs__buff_2 hold198 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[49][1] ),
    .Y(net363));
 sky130_as_sc_hs__buff_2 hold199 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[20][1] ),
    .Y(net364));
 sky130_as_sc_hs__buff_2 hold200 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[51][5] ),
    .Y(net365));
 sky130_as_sc_hs__buff_2 hold201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[29][1] ),
    .Y(net366));
 sky130_as_sc_hs__buff_2 hold202 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_MAR[1] ),
    .Y(net367));
 sky130_as_sc_hs__buff_2 hold203 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[25][2] ),
    .Y(net368));
 sky130_as_sc_hs__buff_2 hold204 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[48][3] ),
    .Y(net369));
 sky130_as_sc_hs__buff_2 hold205 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[8][3] ),
    .Y(net370));
 sky130_as_sc_hs__buff_2 hold206 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[8][1] ),
    .Y(net371));
 sky130_as_sc_hs__buff_2 hold207 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[10][5] ),
    .Y(net372));
 sky130_as_sc_hs__buff_2 hold208 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[32][0] ),
    .Y(net373));
 sky130_as_sc_hs__buff_2 hold209 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[9][0] ),
    .Y(net374));
 sky130_as_sc_hs__buff_2 hold210 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[61][5] ),
    .Y(net375));
 sky130_as_sc_hs__buff_2 hold211 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[51][0] ),
    .Y(net376));
 sky130_as_sc_hs__buff_2 hold212 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[27][3] ),
    .Y(net377));
 sky130_as_sc_hs__buff_2 hold213 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[21][1] ),
    .Y(net378));
 sky130_as_sc_hs__buff_2 hold214 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[48][5] ),
    .Y(net379));
 sky130_as_sc_hs__buff_2 hold215 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[52][1] ),
    .Y(net380));
 sky130_as_sc_hs__buff_2 hold216 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[36][2] ),
    .Y(net381));
 sky130_as_sc_hs__buff_2 hold217 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[18][5] ),
    .Y(net382));
 sky130_as_sc_hs__buff_2 hold218 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[21][5] ),
    .Y(net383));
 sky130_as_sc_hs__buff_2 hold219 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[12][2] ),
    .Y(net384));
 sky130_as_sc_hs__buff_2 hold220 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[10][1] ),
    .Y(net385));
 sky130_as_sc_hs__buff_2 hold221 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[28][5] ),
    .Y(net386));
 sky130_as_sc_hs__buff_2 hold222 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[14][1] ),
    .Y(net387));
 sky130_as_sc_hs__buff_2 hold223 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[51][2] ),
    .Y(net388));
 sky130_as_sc_hs__buff_2 hold224 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[35][3] ),
    .Y(net389));
 sky130_as_sc_hs__buff_2 hold225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[34][1] ),
    .Y(net390));
 sky130_as_sc_hs__buff_2 hold226 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[0][3] ),
    .Y(net391));
 sky130_as_sc_hs__buff_2 hold227 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_P[1] ),
    .Y(net392));
 sky130_as_sc_hs__buff_2 hold228 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[5][1] ),
    .Y(net393));
 sky130_as_sc_hs__buff_2 hold229 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[54][5] ),
    .Y(net394));
 sky130_as_sc_hs__buff_2 hold230 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[22][5] ),
    .Y(net395));
 sky130_as_sc_hs__buff_2 hold231 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[10][4] ),
    .Y(net396));
 sky130_as_sc_hs__buff_2 hold232 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[29][5] ),
    .Y(net397));
 sky130_as_sc_hs__buff_2 hold233 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[0][2] ),
    .Y(net398));
 sky130_as_sc_hs__buff_2 hold234 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[17][1] ),
    .Y(net399));
 sky130_as_sc_hs__buff_2 hold235 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[22][2] ),
    .Y(net400));
 sky130_as_sc_hs__buff_2 hold236 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[25][4] ),
    .Y(net401));
 sky130_as_sc_hs__buff_2 hold237 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[56][5] ),
    .Y(net402));
 sky130_as_sc_hs__buff_2 hold238 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[28][3] ),
    .Y(net403));
 sky130_as_sc_hs__buff_2 hold239 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[57][2] ),
    .Y(net404));
 sky130_as_sc_hs__buff_2 hold240 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[2][1] ),
    .Y(net405));
 sky130_as_sc_hs__buff_2 hold241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[0] ),
    .Y(net406));
 sky130_as_sc_hs__buff_2 hold242 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2315_),
    .Y(net407));
 sky130_as_sc_hs__buff_2 hold243 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[6][2] ),
    .Y(net408));
 sky130_as_sc_hs__buff_2 hold244 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[26][1] ),
    .Y(net409));
 sky130_as_sc_hs__buff_2 hold245 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[27][5] ),
    .Y(net410));
 sky130_as_sc_hs__buff_2 hold246 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[55][3] ),
    .Y(net411));
 sky130_as_sc_hs__buff_2 hold247 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[24][4] ),
    .Y(net412));
 sky130_as_sc_hs__buff_2 hold248 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[13][3] ),
    .Y(net413));
 sky130_as_sc_hs__buff_2 hold249 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[55][5] ),
    .Y(net414));
 sky130_as_sc_hs__buff_2 hold250 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[13][0] ),
    .Y(net415));
 sky130_as_sc_hs__buff_2 hold251 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[61][0] ),
    .Y(net416));
 sky130_as_sc_hs__buff_2 hold252 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[4] ),
    .Y(net417));
 sky130_as_sc_hs__buff_2 hold253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[6][4] ),
    .Y(net418));
 sky130_as_sc_hs__buff_2 hold254 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[47][1] ),
    .Y(net419));
 sky130_as_sc_hs__buff_2 hold255 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[50][0] ),
    .Y(net420));
 sky130_as_sc_hs__buff_2 hold256 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[61][4] ),
    .Y(net421));
 sky130_as_sc_hs__buff_2 hold257 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[39][2] ),
    .Y(net422));
 sky130_as_sc_hs__buff_2 hold258 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[43][3] ),
    .Y(net423));
 sky130_as_sc_hs__buff_2 hold259 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[46][0] ),
    .Y(net424));
 sky130_as_sc_hs__buff_2 hold260 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[24][5] ),
    .Y(net425));
 sky130_as_sc_hs__buff_2 hold261 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[19][5] ),
    .Y(net426));
 sky130_as_sc_hs__buff_2 hold262 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[45][4] ),
    .Y(net427));
 sky130_as_sc_hs__buff_2 hold263 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[36][4] ),
    .Y(net428));
 sky130_as_sc_hs__buff_2 hold264 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[26][4] ),
    .Y(net429));
 sky130_as_sc_hs__buff_2 hold265 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[12][0] ),
    .Y(net430));
 sky130_as_sc_hs__buff_2 hold266 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[24][1] ),
    .Y(net431));
 sky130_as_sc_hs__buff_2 hold267 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[14][4] ),
    .Y(net432));
 sky130_as_sc_hs__buff_2 hold268 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[56][4] ),
    .Y(net433));
 sky130_as_sc_hs__buff_2 hold269 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[9][5] ),
    .Y(net434));
 sky130_as_sc_hs__buff_2 hold270 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[23][3] ),
    .Y(net435));
 sky130_as_sc_hs__buff_2 hold271 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[49][4] ),
    .Y(net436));
 sky130_as_sc_hs__buff_2 hold272 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[0][5] ),
    .Y(net437));
 sky130_as_sc_hs__buff_2 hold273 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[31][2] ),
    .Y(net438));
 sky130_as_sc_hs__buff_2 hold274 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[55][4] ),
    .Y(net439));
 sky130_as_sc_hs__buff_2 hold275 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[20][2] ),
    .Y(net440));
 sky130_as_sc_hs__buff_2 hold276 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[2][3] ),
    .Y(net441));
 sky130_as_sc_hs__buff_2 hold277 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[34][2] ),
    .Y(net442));
 sky130_as_sc_hs__buff_2 hold278 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_MAR[0] ),
    .Y(net443));
 sky130_as_sc_hs__buff_2 hold279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[16][5] ),
    .Y(net444));
 sky130_as_sc_hs__buff_2 hold280 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[13][1] ),
    .Y(net445));
 sky130_as_sc_hs__buff_2 hold281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[2][4] ),
    .Y(net446));
 sky130_as_sc_hs__buff_2 hold282 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[33][3] ),
    .Y(net447));
 sky130_as_sc_hs__buff_2 hold283 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_B[4] ),
    .Y(net448));
 sky130_as_sc_hs__buff_2 hold284 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2342_),
    .Y(net449));
 sky130_as_sc_hs__buff_2 hold285 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[50][1] ),
    .Y(net450));
 sky130_as_sc_hs__buff_2 hold286 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[19][0] ),
    .Y(net451));
 sky130_as_sc_hs__buff_2 hold287 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[61][2] ),
    .Y(net452));
 sky130_as_sc_hs__buff_2 hold288 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[16][2] ),
    .Y(net453));
 sky130_as_sc_hs__buff_2 hold289 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[24][2] ),
    .Y(net454));
 sky130_as_sc_hs__buff_2 hold290 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[47][4] ),
    .Y(net455));
 sky130_as_sc_hs__buff_2 hold291 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[8][4] ),
    .Y(net456));
 sky130_as_sc_hs__buff_2 hold292 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[0][4] ),
    .Y(net457));
 sky130_as_sc_hs__buff_2 hold293 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[4][4] ),
    .Y(net458));
 sky130_as_sc_hs__buff_2 hold294 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[4][2] ),
    .Y(net459));
 sky130_as_sc_hs__buff_2 hold295 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[1] ),
    .Y(net460));
 sky130_as_sc_hs__buff_2 hold296 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2316_),
    .Y(net461));
 sky130_as_sc_hs__buff_2 hold297 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[22][0] ),
    .Y(net462));
 sky130_as_sc_hs__buff_2 hold298 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[10][3] ),
    .Y(net463));
 sky130_as_sc_hs__buff_2 hold299 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[1][1] ),
    .Y(net464));
 sky130_as_sc_hs__buff_2 hold300 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[16][3] ),
    .Y(net465));
 sky130_as_sc_hs__buff_2 hold301 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[37][3] ),
    .Y(net466));
 sky130_as_sc_hs__buff_2 hold302 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[7][1] ),
    .Y(net467));
 sky130_as_sc_hs__buff_2 hold303 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[49][3] ),
    .Y(net468));
 sky130_as_sc_hs__buff_2 hold304 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[22][4] ),
    .Y(net469));
 sky130_as_sc_hs__buff_2 hold305 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[1][0] ),
    .Y(net470));
 sky130_as_sc_hs__buff_2 hold306 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[29][4] ),
    .Y(net471));
 sky130_as_sc_hs__buff_2 hold307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[3][3] ),
    .Y(net472));
 sky130_as_sc_hs__buff_2 hold308 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[5][0] ),
    .Y(net473));
 sky130_as_sc_hs__buff_2 hold309 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[52][3] ),
    .Y(net474));
 sky130_as_sc_hs__buff_2 hold310 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[42][0] ),
    .Y(net475));
 sky130_as_sc_hs__buff_2 hold311 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[35][5] ),
    .Y(net476));
 sky130_as_sc_hs__buff_2 hold312 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[0][0] ),
    .Y(net477));
 sky130_as_sc_hs__buff_2 hold313 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[17][5] ),
    .Y(net478));
 sky130_as_sc_hs__buff_2 hold314 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[42][3] ),
    .Y(net479));
 sky130_as_sc_hs__buff_2 hold315 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[8][2] ),
    .Y(net480));
 sky130_as_sc_hs__buff_2 hold316 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[29][2] ),
    .Y(net481));
 sky130_as_sc_hs__buff_2 hold317 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[6][5] ),
    .Y(net482));
 sky130_as_sc_hs__buff_2 hold318 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[25][3] ),
    .Y(net483));
 sky130_as_sc_hs__buff_2 hold319 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[41][3] ),
    .Y(net484));
 sky130_as_sc_hs__buff_2 hold320 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[32][1] ),
    .Y(net485));
 sky130_as_sc_hs__buff_2 hold321 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[1][5] ),
    .Y(net486));
 sky130_as_sc_hs__buff_2 hold322 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[47][3] ),
    .Y(net487));
 sky130_as_sc_hs__buff_2 hold323 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[51][1] ),
    .Y(net488));
 sky130_as_sc_hs__buff_2 hold324 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[51][4] ),
    .Y(net489));
 sky130_as_sc_hs__buff_2 hold325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[21][2] ),
    .Y(net490));
 sky130_as_sc_hs__buff_2 hold326 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[13][5] ),
    .Y(net491));
 sky130_as_sc_hs__buff_2 hold327 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[5][3] ),
    .Y(net492));
 sky130_as_sc_hs__buff_2 hold328 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[23][1] ),
    .Y(net493));
 sky130_as_sc_hs__buff_2 hold329 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[43][4] ),
    .Y(net494));
 sky130_as_sc_hs__buff_2 hold330 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[50][5] ),
    .Y(net495));
 sky130_as_sc_hs__buff_2 hold331 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[34][4] ),
    .Y(net496));
 sky130_as_sc_hs__buff_2 hold332 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[38][0] ),
    .Y(net497));
 sky130_as_sc_hs__buff_2 hold333 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[47][5] ),
    .Y(net498));
 sky130_as_sc_hs__buff_2 hold334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[14][2] ),
    .Y(net499));
 sky130_as_sc_hs__buff_2 hold335 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_B[1] ),
    .Y(net500));
 sky130_as_sc_hs__buff_2 hold336 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2339_),
    .Y(net501));
 sky130_as_sc_hs__buff_2 hold337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[5][4] ),
    .Y(net502));
 sky130_as_sc_hs__buff_2 hold338 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[11][1] ),
    .Y(net503));
 sky130_as_sc_hs__buff_2 hold339 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[18][2] ),
    .Y(net504));
 sky130_as_sc_hs__buff_2 hold340 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[45][2] ),
    .Y(net505));
 sky130_as_sc_hs__buff_2 hold341 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[19][2] ),
    .Y(net506));
 sky130_as_sc_hs__buff_2 hold342 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[38][4] ),
    .Y(net507));
 sky130_as_sc_hs__buff_2 hold343 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[50][2] ),
    .Y(net508));
 sky130_as_sc_hs__buff_2 hold344 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[9][3] ),
    .Y(net509));
 sky130_as_sc_hs__buff_2 hold345 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[38][1] ),
    .Y(net510));
 sky130_as_sc_hs__buff_2 hold346 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[34][5] ),
    .Y(net511));
 sky130_as_sc_hs__buff_2 hold347 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[2][2] ),
    .Y(net512));
 sky130_as_sc_hs__buff_2 hold348 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[32][5] ),
    .Y(net513));
 sky130_as_sc_hs__buff_2 hold349 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[55][2] ),
    .Y(net514));
 sky130_as_sc_hs__buff_2 hold350 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[54][4] ),
    .Y(net515));
 sky130_as_sc_hs__buff_2 hold351 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[39][3] ),
    .Y(net516));
 sky130_as_sc_hs__buff_2 hold352 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[53][2] ),
    .Y(net517));
 sky130_as_sc_hs__buff_2 hold353 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[43][5] ),
    .Y(net518));
 sky130_as_sc_hs__buff_2 hold354 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[18][3] ),
    .Y(net519));
 sky130_as_sc_hs__buff_2 hold355 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[7][4] ),
    .Y(net520));
 sky130_as_sc_hs__buff_2 hold356 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[62][3] ),
    .Y(net521));
 sky130_as_sc_hs__buff_2 hold357 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[41][1] ),
    .Y(net522));
 sky130_as_sc_hs__buff_2 hold358 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[8][5] ),
    .Y(net523));
 sky130_as_sc_hs__buff_2 hold359 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[42][1] ),
    .Y(net524));
 sky130_as_sc_hs__buff_2 hold360 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[49][5] ),
    .Y(net525));
 sky130_as_sc_hs__buff_2 hold361 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[48][4] ),
    .Y(net526));
 sky130_as_sc_hs__buff_2 hold362 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[29][0] ),
    .Y(net527));
 sky130_as_sc_hs__buff_2 hold363 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[56][2] ),
    .Y(net528));
 sky130_as_sc_hs__buff_2 hold364 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[15][1] ),
    .Y(net529));
 sky130_as_sc_hs__buff_2 hold365 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[31][5] ),
    .Y(net530));
 sky130_as_sc_hs__buff_2 hold366 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[7][3] ),
    .Y(net531));
 sky130_as_sc_hs__buff_2 hold367 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[56][0] ),
    .Y(net532));
 sky130_as_sc_hs__buff_2 hold368 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_B[0] ),
    .Y(net533));
 sky130_as_sc_hs__buff_2 hold369 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2337_),
    .Y(net534));
 sky130_as_sc_hs__buff_2 hold370 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[30][3] ),
    .Y(net535));
 sky130_as_sc_hs__buff_2 hold371 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[32][4] ),
    .Y(net536));
 sky130_as_sc_hs__buff_2 hold372 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[53][4] ),
    .Y(net537));
 sky130_as_sc_hs__buff_2 hold373 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[42][2] ),
    .Y(net538));
 sky130_as_sc_hs__buff_2 hold374 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[50][3] ),
    .Y(net539));
 sky130_as_sc_hs__buff_2 hold375 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[46][3] ),
    .Y(net540));
 sky130_as_sc_hs__buff_2 hold376 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[38][3] ),
    .Y(net541));
 sky130_as_sc_hs__buff_2 hold377 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[26][2] ),
    .Y(net542));
 sky130_as_sc_hs__buff_2 hold378 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[5][5] ),
    .Y(net543));
 sky130_as_sc_hs__buff_2 hold379 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[23][2] ),
    .Y(net544));
 sky130_as_sc_hs__buff_2 hold380 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[52][5] ),
    .Y(net545));
 sky130_as_sc_hs__buff_2 hold381 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[53][5] ),
    .Y(net546));
 sky130_as_sc_hs__buff_2 hold382 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[46][5] ),
    .Y(net547));
 sky130_as_sc_hs__buff_2 hold383 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[36][3] ),
    .Y(net548));
 sky130_as_sc_hs__buff_2 hold384 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[7][0] ),
    .Y(net549));
 sky130_as_sc_hs__buff_2 hold385 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[11][5] ),
    .Y(net550));
 sky130_as_sc_hs__buff_2 hold386 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[3][0] ),
    .Y(net551));
 sky130_as_sc_hs__buff_2 hold387 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[50][4] ),
    .Y(net552));
 sky130_as_sc_hs__buff_2 hold388 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[44][5] ),
    .Y(net553));
 sky130_as_sc_hs__buff_2 hold389 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[41][0] ),
    .Y(net554));
 sky130_as_sc_hs__buff_2 hold390 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[30][5] ),
    .Y(net555));
 sky130_as_sc_hs__buff_2 hold391 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_flags[1] ),
    .Y(net556));
 sky130_as_sc_hs__buff_2 hold392 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[18][4] ),
    .Y(net557));
 sky130_as_sc_hs__buff_2 hold393 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[29][3] ),
    .Y(net558));
 sky130_as_sc_hs__buff_2 hold394 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[16][4] ),
    .Y(net559));
 sky130_as_sc_hs__buff_2 hold395 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_A[0] ),
    .Y(net560));
 sky130_as_sc_hs__buff_2 hold396 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[9][1] ),
    .Y(net561));
 sky130_as_sc_hs__buff_2 hold397 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[3][1] ),
    .Y(net562));
 sky130_as_sc_hs__buff_2 hold398 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[1][2] ),
    .Y(net563));
 sky130_as_sc_hs__buff_2 hold399 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_flags[0] ),
    .Y(net564));
 sky130_as_sc_hs__buff_2 hold400 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[45][5] ),
    .Y(net565));
 sky130_as_sc_hs__buff_2 hold401 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_A[3] ),
    .Y(net566));
 sky130_as_sc_hs__buff_2 hold402 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[41][2] ),
    .Y(net567));
 sky130_as_sc_hs__buff_2 hold403 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[17][4] ),
    .Y(net568));
 sky130_as_sc_hs__buff_2 hold404 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[1][3] ),
    .Y(net569));
 sky130_as_sc_hs__buff_2 hold405 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_A[5] ),
    .Y(net570));
 sky130_as_sc_hs__buff_2 hold406 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\ROM_spi_cycle[4] ),
    .Y(net571));
 sky130_as_sc_hs__buff_2 hold407 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[8][0] ),
    .Y(net572));
 sky130_as_sc_hs__buff_2 hold408 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[62][5] ),
    .Y(net573));
 sky130_as_sc_hs__buff_2 hold409 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_PC[3] ),
    .Y(net574));
 sky130_as_sc_hs__buff_2 hold410 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(_2318_),
    .Y(net575));
 sky130_as_sc_hs__buff_2 hold411 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[2][5] ),
    .Y(net576));
 sky130_as_sc_hs__buff_2 hold412 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\ROM_spi_cycle[2] ),
    .Y(net577));
 sky130_as_sc_hs__buff_2 hold413 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[44][4] ),
    .Y(net578));
 sky130_as_sc_hs__buff_2 hold414 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\imm_buff[5] ),
    .Y(net579));
 sky130_as_sc_hs__buff_2 hold415 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[62][4] ),
    .Y(net580));
 sky130_as_sc_hs__buff_2 hold416 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[62][1] ),
    .Y(net581));
 sky130_as_sc_hs__buff_2 hold417 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\last_A[4] ),
    .Y(net582));
 sky130_as_sc_hs__buff_2 hold418 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[28][4] ),
    .Y(net583));
 sky130_as_sc_hs__buff_2 hold419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(compat),
    .Y(net584));
 sky130_as_sc_hs__buff_2 hold420 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[19][4] ),
    .Y(net585));
 sky130_as_sc_hs__buff_2 hold421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\ROM_spi_cycle[1] ),
    .Y(net586));
 sky130_as_sc_hs__buff_2 hold422 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[62][2] ),
    .Y(net587));
 sky130_as_sc_hs__buff_2 hold423 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\RAM[23][4] ),
    .Y(net588));
 sky130_as_sc_hs__buff_2 hold424 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\imm_buff[3] ),
    .Y(net589));
 sky130_as_sc_hs__buff_2 hold425 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\instr_cycle[1] ),
    .Y(net590));
 sky130_as_sc_hs__buff_2 hold426 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\imm_buff[4] ),
    .Y(net591));
 sky130_as_sc_hs__buff_2 hold427 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\PC[5] ),
    .Y(net592));
 sky130_as_sc_hs__buff_2 hold428 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\ROM_addr_buff[2] ),
    .Y(net593));
 sky130_as_sc_hs__buff_2 hold429 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND),
    .VNB(VGND),
    .A(\instr_cycle[1] ),
    .Y(net594));
 sky130_as_sc_hs__decap_16 FILLER_0_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_0_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_0_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_45 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_73 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_129 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_157 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_185 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_213 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_269 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_297 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_353 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_381 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_409 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_437 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_465 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_493 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_521 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_549 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_577 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_605 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_633 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_661 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_0_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_0_689 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_0_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_0_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_0_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_1_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_353 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_369 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_385 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_425 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_441 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_465 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_1_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_1_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_1_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_1_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_1_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_2_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_2_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_325 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_341 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_357 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_381 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_397 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_413 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_437 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_453 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_469 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_509 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_525 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_2_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_2_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_2_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_2_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_2_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_3_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_353 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_369 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_385 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_425 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_441 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_465 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_3_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_3_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_3_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_3_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_3_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_4_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_4_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_325 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_341 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_357 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_381 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_397 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_413 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_437 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_453 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_469 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_509 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_525 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_4_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_4_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_4_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_4_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_4_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_5_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_353 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_369 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_385 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_425 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_441 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_465 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_5_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_5_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_5_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_5_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_5_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_6_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_6_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_325 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_341 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_357 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_381 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_397 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_413 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_437 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_453 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_469 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_509 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_525 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_6_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_6_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_6_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_6_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_6_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_7_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_353 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_369 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_385 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_425 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_441 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_465 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_7_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_7_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_7_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_7_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_7_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_8_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_8_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_173 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_269 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_285 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_325 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_341 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_357 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_381 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_397 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_413 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_437 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_453 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_469 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_509 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_525 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_8_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_8_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_8_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_8_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_8_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_9_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_73 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_185 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_268 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_272 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_9_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_297 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_353 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_369 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_385 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_425 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_441 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_465 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_9_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_9_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_9_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_9_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_9_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_10_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_10_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_29 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_77 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_101 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_117 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_135 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_10_139 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_10_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_153 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_10_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_10_213 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_221 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_225 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_10_232 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_10_240 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_10_267 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_287 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_303 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_10_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_10_309 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_317 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_335 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_10_339 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_344 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_360 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_381 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_397 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_413 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_437 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_453 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_469 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_509 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_525 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_10_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_10_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_10_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_10_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_10_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_11_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_11_73 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_81 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_11_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_11_105 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_11_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_132 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_11_139 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_11_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_11_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_11_207 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_11_212 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_220 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_273 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_11_295 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_11_300 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_308 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_11_312 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_366 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_11_382 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_11_390 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_425 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_441 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_11_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_465 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_11_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_11_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_11_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_11_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_11_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_11_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_11_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_11_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_12_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_12_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_12_29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_35 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_12_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_12_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_12_115 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_12_135 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_141 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_12_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_12_208 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_12_250 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_257 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_12_309 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_369 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_385 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_401 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_437 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_453 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_469 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_509 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_525 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_12_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_12_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_12_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_12_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_12_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_13_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_13_45 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_13_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_13_88 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_13_103 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_13_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_129 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_13_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_13_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_13_180 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_210 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_13_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_13_265 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_13_291 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_13_316 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_332 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_13_351 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_385 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_425 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_441 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_465 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_13_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_13_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_13_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_13_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_13_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_14_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_14_52 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_14_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_99 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_14_107 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_14_139 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_14_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_14_149 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_160 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_14_180 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_14_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_217 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_14_221 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_257 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_14_270 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_278 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_14_296 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_14_343 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_351 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_14_355 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_392 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_14_408 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_416 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_14_421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_427 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_443 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_459 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_14_475 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_509 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_525 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_14_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_14_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_14_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_14_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_14_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_14_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_14_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_15_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_15_11 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_15_54 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_92 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_142 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_15_146 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_161 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_15_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_177 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_15_205 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_213 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_217 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_15_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_15_249 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_15_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_289 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_15_293 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_15_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_345 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_15_358 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_366 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_15_379 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_387 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_15_391 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_397 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_15_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_15_457 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_467 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_15_483 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_15_503 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_15_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_15_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_15_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_15_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_15_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_15_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_15_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_3 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_16_29 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_16_52 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_16_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_16_89 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_16_104 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_16_129 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_16_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_170 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_174 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_16_216 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_16_240 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_16_250 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_16_257 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_16_268 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_16_292 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_16_319 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_16_336 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_369 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_16_376 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_16_454 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_16_475 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_477 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_16_522 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_16_530 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_16_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_16_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_16_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_16_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_16_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_16_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_17_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_17_43 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_17_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_65 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_17_69 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_90 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_17_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_17_127 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_17_149 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_188 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_17_203 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_17_215 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_223 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_17_229 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_17_259 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_263 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_268 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_300 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_316 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_321 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_348 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_387 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_17_426 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_17_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_17_496 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_529 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_17_545 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_17_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_17_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_17_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_17_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_17_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_17_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_17_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_17_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_17_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_18_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_18_39 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_18_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_63 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_67 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_18_89 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_111 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_18_127 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_18_135 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_141 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_18_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_18_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_18_221 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_263 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_18_300 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_18_328 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_18_336 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_18_362 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_18_379 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_18_384 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_18_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_421 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_18_428 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_18_455 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_18_524 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_18_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_18_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_18_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_18_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_18_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_18_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_7 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_19_33 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_19_54 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_19_67 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_19_79 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_105 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_19_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_117 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_19_140 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_151 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_19_163 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_19_167 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_19_187 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_19_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_19_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_19_233 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_19_249 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_19_264 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_272 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_19_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_286 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_19_298 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_19_311 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_337 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_19_363 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_19_367 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_378 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_382 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_19_393 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_19_408 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_414 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_430 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_434 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_19_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_19_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_457 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_461 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_19_474 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_482 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_19_528 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_544 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_19_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_19_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_19_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_19_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_19_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_19_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_20_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_20_60 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_20_83 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_108 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_112 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_20_138 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_20_145 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_20_153 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_20_187 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_20_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_201 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_20_237 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_20_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_20_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_20_264 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_272 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_20_294 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_20_309 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_20_329 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_20_349 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_20_365 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_373 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_20_405 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_413 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_20_425 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_20_429 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_450 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_20_466 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_20_474 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_20_477 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_20_520 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_528 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_20_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_20_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_20_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_20_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_20_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_20_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_21_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_21_11 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_27 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_21_34 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_38 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_21_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_65 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_21_69 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_21_75 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_146 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_21_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_183 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_21_193 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_201 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_235 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_21_257 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_331 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_335 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_361 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_21_365 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_375 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_21_379 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_21_390 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_403 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_408 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_21_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_21_457 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_488 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_21_492 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_528 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_544 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_21_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_21_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_21_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_21_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_21_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_21_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_3 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_22_25 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_22_49 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_22_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_89 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_22_105 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_117 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_22_139 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_22_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_22_194 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_22_201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_22_242 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_22_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_265 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_22_297 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_22_323 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_22_331 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_360 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_22_369 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_22_408 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_22_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_431 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_22_491 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_22_524 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_22_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_22_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_22_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_22_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_22_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_22_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_23_30 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_23_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_23_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_70 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_23_83 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_23_95 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_23_101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_23_123 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_23_143 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_169 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_23_205 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_23_213 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_239 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_23_243 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_23_285 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_23_360 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_23_403 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_23_407 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_432 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_23_446 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_23_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_457 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_483 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_487 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_23_509 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_23_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_23_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_23_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_23_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_23_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_23_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_23_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_7 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_24_29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_24_34 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_65 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_24_83 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_24_104 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_24_128 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_136 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_24_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_159 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_24_163 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_24_175 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_24_201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_212 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_228 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_24_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_24_267 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_283 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_299 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_24_303 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_319 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_24_355 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_24_363 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_24_365 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_411 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_24_415 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_435 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_24_443 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_24_448 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_24_464 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_472 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_24_497 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_528 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_24_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_24_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_24_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_24_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_24_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_24_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_25_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_15 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_25_22 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_52 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_25_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_65 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_69 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_25_99 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_103 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_25_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_25_156 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_173 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_208 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_25_229 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_25_261 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_265 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_281 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_25_288 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_296 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_300 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_311 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_322 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_25_327 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_335 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_341 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_346 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_357 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_25_368 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_384 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_25_391 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_25_393 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_401 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_406 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_417 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_433 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_437 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_468 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_472 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_497 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_25_505 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_535 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_25_551 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_25_559 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_25_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_25_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_25_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_25_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_25_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_25_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_3 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_26_25 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_26_33 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_26_73 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_26_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_26_99 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_123 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_26_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_26_194 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_26_210 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_221 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_26_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_26_250 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_286 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_26_338 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_26_369 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_377 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_26_381 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_26_405 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_429 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_433 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_26_465 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_26_496 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_26_530 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_26_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_26_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_26_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_26_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_26_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_26_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_27_3 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_27_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_71 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_75 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_167 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_175 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_27_212 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_220 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_235 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_335 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_27_342 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_27_368 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_376 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_391 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_27_403 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_27_470 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_27_505 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_536 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_27_552 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_27_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_27_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_27_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_27_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_27_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_27_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_27_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_7 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_28_33 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_28_56 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_28_72 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_28_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_28_115 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_126 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_130 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_28_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_28_160 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_28_179 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_197 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_28_212 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_28_220 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_28_232 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_28_240 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_28_294 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_28_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_28_309 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_28_324 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_338 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_28_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_28_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_28_407 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_28_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_28_427 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_435 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_443 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_28_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_28_497 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_28_512 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_28_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_28_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_28_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_28_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_28_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_28_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_19 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_29_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_29_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_65 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_69 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_29_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_113 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_29_156 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_29_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_29_222 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_233 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_247 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_29_290 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_298 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_29_328 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_29_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_345 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_350 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_354 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_29_364 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_372 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_376 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_29_386 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_29_401 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_29_409 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_415 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_29_420 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_29_428 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_449 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_29_471 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_29_488 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_505 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_29_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_29_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_29_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_29_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_29_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_29_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_29_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_29_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_30_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_15 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_30_33 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_52 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_30_68 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_30_115 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_30_155 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_176 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_30_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_30_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_201 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_30_233 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_30_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_259 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_30_282 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_30_309 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_325 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_341 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_30_345 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_385 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_30_401 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_30_413 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_30_418 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_30_465 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_477 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_30_494 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_502 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_30_506 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_30_531 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_30_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_30_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_30_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_30_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_30_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_30_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_7 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_31_49 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_31_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_107 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_31_111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_31_117 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_31_157 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_31_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_31_198 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_206 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_31_223 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_31_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_233 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_31_237 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_31_285 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_31_293 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_31_334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_31_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_31_397 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_31_443 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_468 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_31_500 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_31_505 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_513 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_535 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_31_551 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_31_559 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_31_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_31_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_31_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_31_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_31_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_31_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_32_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_32_29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_32_35 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_32_56 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_32_64 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_32_79 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_85 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_32_98 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_114 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_32_151 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_32_159 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_32_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_32_201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_212 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_32_235 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_239 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_32_250 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_263 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_280 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_296 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_323 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_327 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_32_353 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_384 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_400 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_404 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_32_411 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_32_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_32_431 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_439 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_32_475 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_504 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_32_508 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_32_530 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_543 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_559 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_32_575 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_583 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_32_587 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_32_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_32_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_32_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_32_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_32_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_33_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_33_32 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_33_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_33_65 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_33_71 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_107 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_33_111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_33_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_121 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_125 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_33_132 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_33_160 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_33_182 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_190 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_33_194 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_33_239 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_247 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_33_278 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_33_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_33_289 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_33_301 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_33_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_33_358 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_375 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_33_379 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_33_403 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_33_436 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_444 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_33_467 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_475 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_33_479 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_505 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_33_518 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_33_558 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_33_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_33_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_33_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_33_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_33_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_33_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_34_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_34_39 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_55 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_34_59 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_80 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_34_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_110 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_126 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_34_173 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_182 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_186 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_34_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_34_207 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_34_219 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_34_224 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_244 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_34_260 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_34_280 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_292 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_34_296 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_34_322 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_34_338 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_350 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_34_354 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_375 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_379 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_34_415 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_34_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_433 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_34_437 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_34_466 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_34_474 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_34_477 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_34_489 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_34_501 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_34_530 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_537 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_545 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_34_577 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_34_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_34_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_34_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_34_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_34_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_34_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_35_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_35_15 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_35_50 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_35_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_35_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_35_119 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_35_179 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_35_215 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_35_223 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_35_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_35_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_35_286 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_35_290 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_35_326 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_35_334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_35_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_35_345 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_35_364 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_383 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_35_391 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_35_393 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_35_401 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_35_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_35_499 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_538 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_554 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_35_558 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_593 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_35_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_35_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_35_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_35_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_35_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_35_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_35_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_36_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_44 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_36_70 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_36_77 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_36_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_114 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_36_118 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_36_155 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_36_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_36_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_36_253 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_36_266 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_36_278 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_36_286 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_36_331 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_335 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_363 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_36_376 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_36_397 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_405 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_435 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_439 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_36_459 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_36_470 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_36_510 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_36_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_549 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_36_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_36_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_621 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_637 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_36_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_36_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_661 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_36_677 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_693 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_36_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_36_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_36_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_37_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_44 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_37_71 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_79 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_83 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_37_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_37_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_121 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_125 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_140 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_37_155 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_163 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_167 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_179 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_194 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_37_205 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_209 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_37_218 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_37_222 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_229 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_244 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_37_248 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_37_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_289 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_37_308 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_37_322 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_37_357 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_364 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_37_390 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_402 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_422 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_443 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_37_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_37_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_455 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_37_459 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_37_549 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_37_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_577 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_37_586 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_37_602 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_610 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_37_614 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_37_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_37_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_37_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_37_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_37_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_38_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_38_54 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_58 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_38_70 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_78 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_96 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_107 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_123 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_127 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_38_141 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_38_162 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_166 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_181 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_227 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_243 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_247 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_276 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_292 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_296 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_302 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_306 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_347 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_358 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_365 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_401 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_38_421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_450 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_454 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_38_481 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_512 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_528 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_38_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_541 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_38_545 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_38_573 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_599 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_615 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_38_631 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_38_645 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_655 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_38_671 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_38_687 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_695 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_38_699 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_38_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_38_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_39_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_39_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_39_15 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_39_42 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_39_67 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_39_83 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_39_91 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_39_106 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_39_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_39_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_39_158 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_39_169 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_39_182 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_39_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_39_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_39_229 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_39_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_39_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_39_285 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_39_331 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_39_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_39_349 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_39_369 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_39_378 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_39_390 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_39_397 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_39_405 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_39_409 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_39_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_39_453 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_39_477 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_39_485 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_39_489 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_39_500 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_39_509 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_39_525 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_39_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_39_558 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_39_589 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_39_597 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_39_604 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_39_612 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_39_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_39_621 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_39_633 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_39_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_39_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_39_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_39_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_39_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_40_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_40_23 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_40_29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_78 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_40_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_40_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_109 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_40_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_40_201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_40_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_40_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_40_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_40_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_278 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_40_282 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_40_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_40_309 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_40_335 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_40_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_40_375 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_40_407 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_40_418 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_40_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_455 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_40_459 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_40_468 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_40_477 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_40_490 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_40_506 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_514 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_40_518 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_40_531 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_40_537 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_40_543 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_40_565 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_40_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_40_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_40_593 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_40_602 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_40_614 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_40_643 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_40_662 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_40_678 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_694 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_40_698 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_40_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_40_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_41_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_15 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_45 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_41_49 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_41_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_41_73 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_108 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_41_113 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_41_126 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_41_156 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_164 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_192 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_213 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_41_238 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_246 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_281 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_41_285 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_41_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_41_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_353 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_41_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_41_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_453 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_482 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_41_490 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_498 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_41_502 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_41_505 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_513 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_41_529 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_41_545 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_553 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_41_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_41_561 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_41_579 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_595 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_41_631 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_41_650 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_41_664 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_41_691 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_41_707 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_41_711 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_42_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_42_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_43 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_42_83 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_42_99 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_42_105 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_42_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_42_117 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_123 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_42_130 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_42_145 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_42_153 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_157 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_42_193 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_42_201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_42_209 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_42_240 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_42_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_42_276 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_280 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_42_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_309 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_42_326 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_42_334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_42_342 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_42_358 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_42_365 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_42_394 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_42_402 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_42_433 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_42_464 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_42_471 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_42_475 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_42_485 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_42_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_42_541 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_42_559 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_42_567 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_42_571 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_42_577 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_42_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_604 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_42_619 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_42_642 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_42_645 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_42_662 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_42_670 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_42_680 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_42_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_42_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_42_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_43_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_43_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_43_37 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_43_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_43_84 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_43_92 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_96 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_43_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_43_129 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_43_133 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_43_165 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_43_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_180 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_43_196 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_43_204 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_43_229 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_43_251 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_43_270 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_278 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_43_302 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_43_307 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_321 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_43_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_43_345 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_43_361 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_43_365 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_43_382 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_390 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_43_393 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_43_401 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_43_405 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_43_418 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_422 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_465 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_43_479 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_43_499 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_43_519 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_535 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_43_559 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_43_561 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_43_583 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_43_591 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_43_610 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_614 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_43_617 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_43_625 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_43_630 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_43_646 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_43_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_43_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_43_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_44_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_44_39 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_47 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_55 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_44_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_44_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_44_93 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_44_117 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_44_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_44_160 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_44_168 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_44_173 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_44_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_44_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_208 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_44_212 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_44_253 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_44_265 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_44_277 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_44_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_44_349 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_357 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_44_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_44_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_44_400 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_44_425 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_465 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_44_474 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_44_477 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_44_482 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_44_498 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_506 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_44_513 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_44_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_44_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_44_537 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_44_554 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_582 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_44_586 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_44_589 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_44_618 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_634 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_679 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_696 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_44_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_44_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_45_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_45_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_45_37 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_45_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_45_88 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_45_96 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_45_104 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_45_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_45_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_45_209 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_45_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_45_271 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_45_275 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_45_313 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_45_335 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_45_343 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_45_351 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_45_393 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_45_405 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_45_420 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_45_428 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_45_432 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_45_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_45_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_45_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_45_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_45_505 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_45_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_45_537 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_45_545 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_45_584 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_45_594 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_45_603 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_45_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_45_625 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_45_666 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_45_670 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_45_688 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_45_704 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_45_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_46_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_46_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_46_29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_46_41 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_46_85 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_46_92 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_46_133 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_46_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_46_162 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_46_206 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_46_210 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_46_263 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_46_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_46_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_46_341 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_46_349 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_46_379 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_46_383 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_46_395 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_46_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_46_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_46_437 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_46_455 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_46_474 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_46_494 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_46_498 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_46_530 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_46_533 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_46_541 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_46_549 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_46_555 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_46_563 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_46_579 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_46_587 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_46_601 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_46_620 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_46_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_46_637 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_46_653 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_46_687 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_46_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_46_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_47_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_47_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_47_15 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_47_50 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_47_54 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_47_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_47_61 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_47_74 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_47_100 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_47_104 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_47_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_47_127 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_47_143 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_47_155 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_163 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_47_174 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_47_195 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_199 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_47_209 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_217 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_47_222 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_47_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_250 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_47_256 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_47_260 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_47_281 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_47_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_47_331 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_335 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_47_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_47_345 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_349 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_47_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_47_423 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_47_427 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_47_440 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_47_459 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_47_497 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_47_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_47_505 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_47_528 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_47_548 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_47_575 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_582 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_47_596 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_47_612 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_47_629 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_47_645 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_47_653 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_657 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_671 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_47_704 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_47_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_48_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_48_29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_48_50 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_62 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_48_114 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_48_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_48_171 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_48_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_205 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_48_209 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_230 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_48_234 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_48_242 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_48_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_48_263 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_48_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_287 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_48_291 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_48_299 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_48_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_48_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_383 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_48_421 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_48_453 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_48_468 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_491 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_48_505 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_48_530 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_48_586 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_48_603 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_48_619 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_48_665 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_680 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_695 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_48_699 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_48_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_48_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_49_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_50 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_54 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_49_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_73 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_88 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_49_103 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_136 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_167 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_203 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_207 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_218 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_251 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_255 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_270 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_274 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_292 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_296 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_49_308 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_49_330 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_49_341 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_49_375 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_391 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_407 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_411 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_446 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_49_453 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_461 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_472 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_49_476 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_49_486 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_490 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_502 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_49_520 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_49_527 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_554 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_558 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_599 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_609 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_49_613 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_49_627 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_49_631 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_49_662 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_670 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_49_685 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_49_708 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_49_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_50_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_50_15 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_50_29 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_50_55 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_50_69 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_80 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_50_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_50_101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_50_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_50_139 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_50_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_50_184 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_50_201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_50_222 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_233 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_50_237 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_50_257 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_50_284 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_333 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_50_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_378 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_50_382 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_50_402 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_50_410 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_50_425 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_50_437 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_50_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_50_457 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_469 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_50_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_50_511 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_528 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_50_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_50_546 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_50_562 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_50_602 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_610 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_50_614 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_50_625 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_50_633 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_50_645 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_50_669 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_50_678 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_50_686 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_50_691 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_50_699 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_50_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_50_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_30 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_68 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_80 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_84 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_99 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_51_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_51_113 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_51_140 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_156 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_164 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_178 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_195 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_199 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_51_222 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_51_240 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_51_288 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_51_305 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_312 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_316 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_51_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_51_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_341 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_377 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_385 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_51_411 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_51_427 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_436 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_444 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_51_464 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_51_487 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_503 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_505 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_516 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_535 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_551 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_559 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_561 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_51_569 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_51_576 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_607 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_624 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_628 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_662 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_51_666 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_51_670 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_51_698 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_51_706 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_51_710 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_52_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_52_63 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_71 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_52_104 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_52_108 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_52_133 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_52_151 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_182 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_52_189 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_52_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_52_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_52_213 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_52_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_52_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_52_296 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_52_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_52_309 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_52_325 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_52_332 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_337 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_52_369 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_52_377 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_381 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_52_413 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_52_421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_52_429 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_52_474 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_489 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_52_507 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_52_515 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_52_526 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_52_552 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_52_568 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_52_576 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_580 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_52_606 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_52_628 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_52_640 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_52_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_52_689 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_52_693 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_52_699 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_52_711 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_53_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_53_7 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_53_34 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_53_42 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_53_50 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_53_54 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_53_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_53_69 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_53_129 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_53_179 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_53_202 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_53_210 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_53_214 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_53_248 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_53_256 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_53_276 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_53_289 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_53_308 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_53_312 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_53_324 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_53_328 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_53_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_53_337 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_53_344 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_53_364 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_53_380 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_53_415 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_53_423 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_53_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_53_456 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_53_479 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_53_497 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_53_543 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_53_550 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_53_558 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_53_561 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_53_569 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_53_612 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_53_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_53_621 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_53_638 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_53_644 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_53_658 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_53_662 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_53_685 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_53_710 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_54_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_54_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_54_29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_54_60 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_54_68 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_54_72 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_54_118 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_54_155 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_54_248 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_54_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_54_261 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_54_269 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_54_306 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_54_317 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_54_349 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_54_358 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_54_365 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_54_374 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_54_382 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_54_418 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_54_421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_54_472 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_54_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_54_481 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_54_519 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_54_524 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_54_533 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_54_542 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_54_550 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_54_554 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_54_578 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_54_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_54_612 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_54_620 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_54_624 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_54_632 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_54_638 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_54_642 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_54_650 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_54_654 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_54_680 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_54_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_54_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_32 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_55_67 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_75 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_55_102 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_55_110 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_55_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_129 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_55_153 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_55_161 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_55_179 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_218 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_55_239 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_55_261 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_266 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_308 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_55_334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_55_351 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_55_373 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_387 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_393 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_55_417 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_425 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_55_449 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_55_458 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_55_466 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_55_482 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_55_493 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_55_512 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_55_528 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_559 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_55_561 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_55_567 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_55_583 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_592 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_55_603 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_55_614 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_55_617 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_55_627 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_55_650 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_55_667 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_55_671 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_55_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_55_689 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_55_710 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_56_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_56_33 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_56_60 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_56_68 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_72 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_83 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_56_91 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_56_95 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_56_108 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_56_116 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_56_129 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_56_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_56_145 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_56_149 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_56_184 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_190 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_56_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_56_301 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_56_305 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_56_309 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_56_322 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_56_357 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_56_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_56_375 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_56_415 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_56_421 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_56_444 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_56_452 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_456 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_477 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_56_513 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_56_521 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_56_525 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_56_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_571 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_587 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_56_602 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_628 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_56_645 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_56_676 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_56_684 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_56_698 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_56_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_57_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_57_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_57_28 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_57_39 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_57_43 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_57_48 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_57_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_57_65 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_57_99 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_57_136 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_57_144 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_57_148 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_57_164 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_57_178 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_57_182 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_57_193 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_57_204 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_57_222 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_57_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_57_250 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_57_273 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_57_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_57_300 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_57_334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_57_351 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_57_413 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_57_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_57_478 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_57_511 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_57_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_57_547 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_57_558 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_57_573 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_57_594 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_57_605 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_57_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_57_627 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_57_660 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_57_684 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_57_710 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_58_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_33 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_58_39 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_58_55 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_59 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_58_91 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_58_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_138 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_58_141 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_58_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_58_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_58_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_264 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_58_290 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_58_298 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_302 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_58_309 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_58_347 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_58_355 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_58_359 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_58_375 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_58_386 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_58_407 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_58_415 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_58_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_58_471 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_493 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_58_514 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_530 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_58_533 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_58_548 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_58_587 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_58_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_593 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_605 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_58_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_58_635 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_58_686 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_58_690 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_58_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_58_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_58_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_59_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_59_44 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_59_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_59_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_84 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_59_97 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_166 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_194 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_59_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_59_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_59_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_59_292 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_59_351 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_375 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_59_415 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_59_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_434 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_446 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_59_461 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_59_469 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_59_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_59_482 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_59_494 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_59_501 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_59_520 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_59_556 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_59_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_638 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_59_643 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_59_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_59_680 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_59_688 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_59_710 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_60_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_60_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_60_29 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_60_65 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_60_69 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_60_89 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_60_105 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_60_112 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_60_120 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_60_139 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_60_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_60_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_60_248 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_60_295 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_60_299 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_60_306 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_60_335 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_60_351 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_60_359 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_60_363 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_60_383 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_60_416 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_60_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_60_425 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_60_450 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_60_454 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_60_475 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_60_491 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_60_507 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_60_515 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_60_548 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_60_556 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_60_589 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_60_631 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_60_645 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_60_651 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_60_659 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_60_663 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_60_690 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_60_698 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_60_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_60_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_61_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_61_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_61_39 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_61_108 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_61_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_61_121 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_61_146 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_61_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_61_194 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_61_206 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_61_222 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_61_234 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_61_255 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_61_271 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_61_297 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_61_341 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_61_353 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_61_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_61_381 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_61_385 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_61_413 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_61_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_61_457 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_61_487 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_61_503 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_61_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_61_509 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_61_516 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_61_525 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_61_550 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_61_588 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_61_596 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_61_608 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_61_636 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_61_652 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_61_660 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_61_671 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_61_673 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_61_704 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_61_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_62_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_62_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_62_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_62_63 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_62_85 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_62_117 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_62_139 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_62_187 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_62_234 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_62_241 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_62_245 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_62_286 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_62_304 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_62_317 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_62_326 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_62_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_62_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_62_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_62_369 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_62_381 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_62_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_62_413 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_62_436 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_62_457 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_62_461 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_62_467 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_62_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_62_485 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_62_517 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_62_525 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_62_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_62_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_62_545 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_62_586 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_62_596 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_62_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_62_645 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_62_653 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_62_683 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_62_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_62_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_62_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_63_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_63_30 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_63_61 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_63_86 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_63_111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_63_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_63_117 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_63_146 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_63_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_63_180 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_63_203 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_63_244 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_63_252 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_63_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_63_299 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_63_319 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_63_327 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_63_331 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_63_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_63_403 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_63_411 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_63_415 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_63_435 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_63_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_63_457 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_63_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_63_485 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_63_527 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_63_543 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_63_559 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_63_561 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_63_567 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_63_575 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_63_582 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_63_608 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_63_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_63_644 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_63_648 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_63_688 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_63_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_64_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_15 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_64_27 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_64_33 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_41 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_64_53 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_64_64 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_64_89 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_64_111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_119 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_123 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_64_129 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_64_147 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_64_178 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_194 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_238 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_242 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_272 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_64_276 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_64_306 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_64_319 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_327 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_64_369 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_64_384 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_64_397 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_413 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_64_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_64_421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_429 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_437 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_64_441 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_64_450 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_64_477 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_485 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_64_497 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_64_526 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_530 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_64_571 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_64_587 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_589 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_64_620 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_628 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_64_634 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_64_642 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_645 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_64_649 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_64_663 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_64_679 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_64_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_64_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_65_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_19 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_65_27 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_65_43 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_65_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_65_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_65_65 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_65_95 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_65_99 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_107 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_65_111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_65_123 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_65_130 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_65_146 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_162 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_65_183 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_191 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_65_225 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_65_241 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_249 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_274 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_278 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_65_281 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_65_326 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_330 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_360 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_368 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_382 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_388 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_65_393 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_65_422 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_65_430 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_446 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_476 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_480 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_502 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_65_536 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_573 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_65_577 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_65_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_65_617 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_625 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_65_629 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_65_635 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_65_678 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_65_708 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_65_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_66_29 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_66_46 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_66_62 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_66_75 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_83 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_66_101 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_66_118 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_139 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_66_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_157 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_161 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_191 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_213 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_238 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_246 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_250 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_253 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_257 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_66_265 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_273 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_277 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_301 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_66_326 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_66_334 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_66_343 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_66_349 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_357 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_388 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_441 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_474 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_66_477 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_66_517 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_525 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_66_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_66_533 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_537 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_571 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_575 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_589 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_66_610 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_66_626 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_642 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_645 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_66_667 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_66_671 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_66_678 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_66_686 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_66_693 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_66_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_66_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_67_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_67_48 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_76 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_152 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_183 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_206 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_210 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_216 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_67_235 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_67_264 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_67_270 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_278 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_67_281 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_67_315 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_67_328 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_67_337 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_67_353 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_361 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_384 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_403 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_67_421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_429 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_67_469 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_67_476 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_484 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_502 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_67_509 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_67_518 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_534 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_67_542 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_570 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_67_587 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_67_602 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_67_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_621 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_629 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_67_645 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_67_686 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_67_690 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_67_710 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_68_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_68_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_68_39 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_68_71 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_68_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_68_124 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_68_141 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_68_145 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_68_182 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_68_207 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_68_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_68_321 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_68_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_68_358 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_68_362 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_68_365 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_68_373 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_68_377 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_68_418 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_68_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_68_425 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_68_445 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_68_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_68_472 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_68_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_68_493 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_68_539 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_68_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_68_589 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_68_620 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_68_628 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_68_633 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_68_695 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_68_699 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_68_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_69_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_69_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_69_46 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_69_50 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_69_61 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_69_87 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_69_105 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_69_123 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_69_127 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_69_136 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_69_144 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_69_174 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_69_185 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_69_193 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_69_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_69_233 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_69_237 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_69_277 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_69_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_69_315 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_69_323 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_69_327 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_69_368 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_69_384 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_69_396 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_69_414 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_69_418 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_69_446 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_69_455 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_69_548 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_69_574 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_69_580 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_69_584 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_69_596 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_69_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_69_632 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_69_654 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_69_684 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_69_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_69_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_70_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_70_11 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_70_47 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_70_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_70_71 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_70_78 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_70_82 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_99 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_70_103 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_70_114 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_130 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_70_134 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_70_145 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_153 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_70_157 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_70_169 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_191 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_70_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_70_201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_70_228 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_236 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_70_240 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_70_263 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_70_288 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_70_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_70_320 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_349 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_70_353 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_70_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_381 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_70_385 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_70_409 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_70_417 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_70_421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_429 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_70_433 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_469 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_70_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_70_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_70_493 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_70_548 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_70_573 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_70_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_70_589 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_70_593 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_70_626 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_70_682 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_70_695 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_70_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_70_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_71_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_71_15 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_71_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_65 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_71_69 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_71_96 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_108 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_118 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_122 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_71_152 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_169 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_173 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_71_189 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_71_235 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_71_251 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_71_267 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_275 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_279 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_71_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_289 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_71_305 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_321 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_325 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_330 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_71_334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_71_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_71_371 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_71_379 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_71_412 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_71_424 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_71_440 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_71_468 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_71_484 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_500 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_71_511 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_71_536 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_552 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_71_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_71_580 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_71_590 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_71_594 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_71_602 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_71_627 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_658 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_671 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_71_678 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_71_687 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_71_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_72_58 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_72_116 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_124 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_163 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_72_167 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_72_197 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_72_229 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_245 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_72_249 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_72_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_259 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_72_266 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_280 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_72_288 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_72_341 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_352 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_362 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_377 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_72_412 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_72_442 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_466 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_487 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_72_491 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_496 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_72_525 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_72_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_72_547 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_567 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_578 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_586 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_72_589 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_628 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_72_632 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_72_643 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_72_645 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_72_658 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_72_666 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_670 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_72_691 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_72_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_72_705 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_73_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_73_53 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_73_111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_73_146 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_73_169 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_73_182 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_73_202 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_73_221 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_73_233 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_73_241 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_73_334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_383 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_410 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_73_414 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_73_439 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_73_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_73_503 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_73_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_73_521 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_527 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_73_531 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_73_543 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_73_551 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_572 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_592 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_600 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_73_604 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_73_611 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_73_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_73_631 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_73_639 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_73_663 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_73_671 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_73_708 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_73_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_74_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_74_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_74_15 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_74_29 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_74_52 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_74_56 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_74_61 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_74_77 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_74_99 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_74_107 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_74_111 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_74_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_74_151 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_74_159 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_74_163 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_74_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_74_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_74_224 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_74_240 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_74_264 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_74_300 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_74_318 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_74_334 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_74_344 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_74_375 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_74_473 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_74_481 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_74_485 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_74_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_74_521 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_74_552 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_74_586 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_74_595 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_74_611 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_74_619 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_74_630 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_74_672 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_74_707 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_74_711 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_75_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_75_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_75_46 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_75_54 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_57 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_75_70 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_86 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_75_93 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_75_101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_75_113 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_75_144 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_75_160 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_169 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_75_176 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_75_192 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_75_200 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_75_204 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_75_235 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_75_262 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_298 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_75_307 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_75_323 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_75_334 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_337 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_75_346 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_75_356 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_75_363 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_75_367 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_371 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_75_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_413 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_75_420 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_75_430 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_75_438 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_75_442 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_75_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_75_461 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_465 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_75_502 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_75_511 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_75_519 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_75_523 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_75_546 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_75_554 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_75_558 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_75_607 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_75_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_75_638 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_75_670 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_75_673 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_75_681 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_75_707 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_75_711 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_76_7 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_76_29 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_76_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_76_85 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_76_97 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_76_124 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_76_137 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_76_151 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_165 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_76_182 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_190 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_76_194 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_76_197 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_76_232 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_248 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_253 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_258 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_264 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_270 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_76_300 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_76_309 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_76_322 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_352 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_407 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_411 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_76_418 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_421 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_76_425 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_76_433 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_76_444 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_460 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_76_464 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_76_472 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_76_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_493 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_505 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_76_519 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_527 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_531 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_76_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_76_541 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_76_550 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_76_557 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_76_573 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_581 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_76_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_76_589 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_76_605 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_76_621 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_629 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_633 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_76_645 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_676 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_76_680 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_76_687 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_76_697 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_76_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_76_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_77_3 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_77_47 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_77_57 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_77_81 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_77_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_77_183 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_77_239 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_77_243 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_77_249 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_77_257 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_77_281 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_77_299 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_77_307 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_77_313 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_77_317 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_77_330 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_77_343 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_77_366 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_77_370 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_77_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_77_406 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_77_410 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_77_442 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_77_449 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_77_453 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_77_479 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_77_515 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_77_529 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_77_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_77_561 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_77_569 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_77_573 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_77_617 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_77_625 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_77_629 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_77_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_77_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_77_710 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_78_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_78_49 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_78_74 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_78_81 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_78_95 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_78_118 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_78_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_78_197 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_78_233 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_78_237 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_78_287 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_78_316 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_78_336 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_78_340 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_78_353 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_78_362 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_78_365 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_78_407 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_78_421 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_78_450 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_78_483 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_78_522 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_78_530 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_78_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_78_559 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_78_623 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_78_712 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_79_3 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_79_11 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_79_15 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_79_51 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_79_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_79_71 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_79_98 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_79_144 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_3 FILLER_79_179 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_79_225 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_79_233 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_79_296 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_79_332 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_79_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_79_363 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_79_379 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_79_387 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_79_391 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_79_393 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_79_401 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_79_445 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_79_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_79_478 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_79_482 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_79_521 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_79_529 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_79_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_79_557 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_79_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_79_615 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_79_617 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_79_625 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_79_629 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_79_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_79_673 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_79_702 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_79_710 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_80_3 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_80_19 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_25 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_80_47 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_55 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_57 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_64 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_80_70 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_80_78 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_80_85 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_101 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_109 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_80_113 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_80_118 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_130 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_80_138 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_141 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_149 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_153 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_80_179 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_195 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_201 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_80_209 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_215 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_225 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_80_259 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_286 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_2 FILLER_80_293 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_80_299 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_309 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_315 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_320 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_329 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_333 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_80_337 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_345 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_349 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_357 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_361 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_80_365 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_381 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_389 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_80_393 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_409 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_419 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_425 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_429 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_4 FILLER_80_443 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_447 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_449 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_457 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_461 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_472 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_80_477 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_493 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_498 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_80_502 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_80_505 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_521 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_529 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_80_533 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_1 FILLER_80_541 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_550 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_80_558 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_80_561 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_577 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_585 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_1 FILLER_80_589 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_602 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_610 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_2 FILLER_80_614 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_16 FILLER_80_617 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_633 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_641 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__decap_16 FILLER_80_649 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_665 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_669 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_80_673 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_681 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_3 FILLER_80_685 (.VNB(VGND),
    .VPB(VPWR),
    .VGND(VGND),
    .VPWR(VPWR));
 sky130_as_sc_hs__fill_8 FILLER_80_692 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__fill_8 FILLER_80_701 (.VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 sky130_as_sc_hs__decap_4 FILLER_80_709 (.VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .VGND(VGND));
 assign uio_oe[6] = net163;
 assign uio_oe[7] = net165;
 assign uio_out[6] = net164;
endmodule
